// Register NVDLA_RBK_S_STATUS_0
#define NVDLA_RBK_S_STATUS_0					32'h11000
#define NVDLA_RBK_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_RBK_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_RBK_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_RBK_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_RBK_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_RBK_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_RBK_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_RBK_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_RBK_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_RBK_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_RBK_S_POINTER_0
#define NVDLA_RBK_S_POINTER_0					32'h11004
#define NVDLA_RBK_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_RBK_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_RBK_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_RBK_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_RBK_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_RBK_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_RBK_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_RBK_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_RBK_D_OP_ENABLE_0
#define NVDLA_RBK_D_OP_ENABLE_0					32'h11008
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_RBK_D_MISC_CFG_0
#define NVDLA_RBK_D_MISC_CFG_0					32'h1100c
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_RANGE			1:0
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_SIZE				2
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_CONTRACT			2'h0
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_SPLIT			2'h1
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_MERGE			2'h2
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_RANGE			9:8
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_FP16			2'h2


// Register NVDLA_RBK_D_DAIN_RAM_TYPE_0
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0					32'h11010
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_RANGE			0:0
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_SIZE				1
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_CVIF			1'h0
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_MCIF			1'h1


// Register NVDLA_RBK_D_DATAIN_SIZE_0_0
#define NVDLA_RBK_D_DATAIN_SIZE_0_0					32'h11014
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_WIDTH_RANGE			12:0
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_WIDTH_SIZE				13
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_HEIGHT_RANGE			28:16
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_HEIGHT_SIZE				13


// Register NVDLA_RBK_D_DATAIN_SIZE_1_0
#define NVDLA_RBK_D_DATAIN_SIZE_1_0					32'h11018
#define NVDLA_RBK_D_DATAIN_SIZE_1_0_DATAIN_CHANNEL_RANGE			12:0
#define NVDLA_RBK_D_DATAIN_SIZE_1_0_DATAIN_CHANNEL_SIZE				13


// Register NVDLA_RBK_D_DAIN_ADDR_HIGH_0
#define NVDLA_RBK_D_DAIN_ADDR_HIGH_0					32'h1101c
#define NVDLA_RBK_D_DAIN_ADDR_HIGH_0_DAIN_ADDR_HIGH_RANGE			31:0
#define NVDLA_RBK_D_DAIN_ADDR_HIGH_0_DAIN_ADDR_HIGH_SIZE				32


// Register NVDLA_RBK_D_DAIN_ADDR_LOW_0
#define NVDLA_RBK_D_DAIN_ADDR_LOW_0					32'h11020
#define NVDLA_RBK_D_DAIN_ADDR_LOW_0_DAIN_ADDR_LOW_RANGE			31:5
#define NVDLA_RBK_D_DAIN_ADDR_LOW_0_DAIN_ADDR_LOW_SIZE				27


// Register NVDLA_RBK_D_DAIN_LINE_STRIDE_0
#define NVDLA_RBK_D_DAIN_LINE_STRIDE_0					32'h11024
#define NVDLA_RBK_D_DAIN_LINE_STRIDE_0_DAIN_LINE_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAIN_LINE_STRIDE_0_DAIN_LINE_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAIN_SURF_STRIDE_0
#define NVDLA_RBK_D_DAIN_SURF_STRIDE_0					32'h11028
#define NVDLA_RBK_D_DAIN_SURF_STRIDE_0_DAIN_SURF_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAIN_SURF_STRIDE_0_DAIN_SURF_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0
#define NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0					32'h1102c
#define NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0_DAIN_PLANAR_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0_DAIN_PLANAR_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAOUT_RAM_TYPE_0
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0					32'h11030
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_RANGE			0:0
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_SIZE				1
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_CVIF			1'h0
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_MCIF			1'h1


// Register NVDLA_RBK_D_DATAOUT_SIZE_1_0
#define NVDLA_RBK_D_DATAOUT_SIZE_1_0					32'h11034
#define NVDLA_RBK_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_RANGE			12:0
#define NVDLA_RBK_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_SIZE				13


// Register NVDLA_RBK_D_DAOUT_ADDR_HIGH_0
#define NVDLA_RBK_D_DAOUT_ADDR_HIGH_0					32'h11038
#define NVDLA_RBK_D_DAOUT_ADDR_HIGH_0_DAOUT_ADDR_HIGH_RANGE			31:0
#define NVDLA_RBK_D_DAOUT_ADDR_HIGH_0_DAOUT_ADDR_HIGH_SIZE				32


// Register NVDLA_RBK_D_DAOUT_ADDR_LOW_0
#define NVDLA_RBK_D_DAOUT_ADDR_LOW_0					32'h1103c
#define NVDLA_RBK_D_DAOUT_ADDR_LOW_0_DAOUT_ADDR_LOW_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_ADDR_LOW_0_DAOUT_ADDR_LOW_SIZE				27


// Register NVDLA_RBK_D_DAOUT_LINE_STRIDE_0
#define NVDLA_RBK_D_DAOUT_LINE_STRIDE_0					32'h11040
#define NVDLA_RBK_D_DAOUT_LINE_STRIDE_0_DAOUT_LINE_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_LINE_STRIDE_0_DAOUT_LINE_STRIDE_SIZE				27


// Register NVDLA_RBK_D_CONTRACT_STRIDE_0_0
#define NVDLA_RBK_D_CONTRACT_STRIDE_0_0					32'h11044
#define NVDLA_RBK_D_CONTRACT_STRIDE_0_0_CONTRACT_STRIDE_0_RANGE			31:5
#define NVDLA_RBK_D_CONTRACT_STRIDE_0_0_CONTRACT_STRIDE_0_SIZE				27


// Register NVDLA_RBK_D_CONTRACT_STRIDE_1_0
#define NVDLA_RBK_D_CONTRACT_STRIDE_1_0					32'h11048
#define NVDLA_RBK_D_CONTRACT_STRIDE_1_0_CONTRACT_STRIDE_1_RANGE			31:5
#define NVDLA_RBK_D_CONTRACT_STRIDE_1_0_CONTRACT_STRIDE_1_SIZE				27


// Register NVDLA_RBK_D_DAOUT_SURF_STRIDE_0
#define NVDLA_RBK_D_DAOUT_SURF_STRIDE_0					32'h1104c
#define NVDLA_RBK_D_DAOUT_SURF_STRIDE_0_DAOUT_SURF_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_SURF_STRIDE_0_DAOUT_SURF_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0
#define NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0					32'h11050
#define NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0_DAOUT_PLANAR_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0_DAOUT_PLANAR_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DECONV_STRIDE_0
#define NVDLA_RBK_D_DECONV_STRIDE_0					32'h11054
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_X_STRIDE_RANGE			4:0
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_X_STRIDE_SIZE				5
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_Y_STRIDE_RANGE			20:16
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_Y_STRIDE_SIZE				5


// Register NVDLA_RBK_D_PERF_ENABLE_0
#define NVDLA_RBK_D_PERF_ENABLE_0					32'h11058
#define NVDLA_RBK_D_PERF_ENABLE_0_PERF_EN_RANGE			0:0
#define NVDLA_RBK_D_PERF_ENABLE_0_PERF_EN_SIZE				1


// Register NVDLA_RBK_D_PERF_READ_STALL_0
#define NVDLA_RBK_D_PERF_READ_STALL_0					32'h1105c
#define NVDLA_RBK_D_PERF_READ_STALL_0_RD_STALL_CNT_RANGE			31:0
#define NVDLA_RBK_D_PERF_READ_STALL_0_RD_STALL_CNT_SIZE				32


// Register NVDLA_RBK_D_PERF_WRITE_STALL_0
#define NVDLA_RBK_D_PERF_WRITE_STALL_0					32'h11060
#define NVDLA_RBK_D_PERF_WRITE_STALL_0_WR_STALL_CNT_RANGE			31:0
#define NVDLA_RBK_D_PERF_WRITE_STALL_0_WR_STALL_CNT_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_RBK	32'h11000
