`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NK6na3mE378GlzxIGWaMd5DMDagwF81guhrTmz37HsTcMhCpKHMHZIa0wIPCmoAuXglaPGtps7LI
ityA46V6tg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D+TO6SfSGUDinzYLaz9SdIF4WhY4zYQQoSYFbZ8fJY9lT56eS1OXtSnZTEy8ELJXRBHOgSorUyus
K5vnayeBS+gjia/mk/M5wMDxLrhhpi5JOcFlEQM03aMdqYM3pQuNR/jsqddSxNwlT04J6vMOG7BO
xtPSdy5In6+3OltlU7E=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQu4CtbDuqvs1PJt8fBD8x3y1o7ApfM7m4TuKWGMHX6g2T0l8f9hLK3eVuUDFWEl3Qa8RX/SedXs
RHTYNsu7LEwtwp5vyH0i5SKvBhqudQon7kKCsiaPVjMJlchpNQyDh8AShPGOfgGRf0NckiS7mnTH
xq0X7n4RTNITGnD48Kukpn54Et+0UARAQi6zNeoLA4W4VAWP4rFTAoHHB3I9wvS9h/cHeaCrmnm/
bPVDxw5FhvHykvzeeurzFp4Qg/iATE7oW4zeao+g2fQPT7mXhpbIvDQoQbidqYzV8uvtprdykYMM
npBXeibmqrdPVdSf0P58VzChnY5sysGzEKYimA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FISISVTuxCDORPkxiQemMoF/Y4djak9O/AftgXIjwVtSRd7vaohVcxXIudX1SdKZKIVYq3zFbqFo
OnxjCnIcJque30/xNbeSFJwzWoEn1/yL8SDx+cNASz9YtTZVcsoLXYzMqlTudu65Qi9kXxtV6kKr
l2s7Oao8wlrnFNwL2KahnqsWa+TD0T/7+wPkWdfz5zbPHmabHHDQOGUhryb7q5tgfEmkULOOIl12
EwXvd+oOeYLPjcuZGzMk7sQX37C4wpAwO1fcKCeaMchWWNoWZjLjSmDbd4fHM7DTxF8VMrXd8SFl
yAEfVIjYwY8Z7A8TvOaXcWWkY3i2/EGDqETLfw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V0DarZWaKeaBKmybJ/G93dmkWSmlFnY/5g+hKP3FuZ8HNasz5GmHJpHG86E/yGJ1wFRigDPTZNXR
xFJFg8H7WgjFXe66yfkLEMusQVwZHaiDgMhrUXBUzEWqTXH83Xde6acKWX9VdjxswHaR9IMWtEPx
aVItmgrmj26PoT0rGEV86iJqQNpwTW0/Xme9O1isHn1rsh7z+P1eu7dhAFi98GBfe6+79LziEsbb
u1Y+zRdAApL2ANkY5yjFRMc2/BSnB1yGM1U5ZfsCYlML41/0CdDx5aI4QPqs+C9iSx7d1iiu3WhN
rChnBdD+wSLPCPU5vTXzRv+c5JV79S0e5394Yg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L/x+xmJXV7qUsSHdMUJn+SI4tfyPZEfZ42z6MDC52y/cMdob46gs3zazJJDwBJln99EpCTqqzyBF
u2Kx7SYDvBYc6xvHT/lXIyDNbI+wh2o/WxeSMEILef0gqFwyW2RtwNppyrQ76GfMaw3HofyR9l7Z
DXW42IjhEaXfLD+RRQI=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B8zopJE9SDlNaEvIu39LxGkQY3MYcfT3GNUdp22wTuy8uuOKZQMWTNM+k+qRco+sDI/8Gwc4b0dE
G7MKERyWv0YyoEjeZPi6MRUoOmFl3gE7R0HWU2V2hjuJP+YaQYj19PmSw1/6HAGN7hfwYTp7UZpa
R4qw/uroN6jDm+NR8AE8kD0xWJkyvDXxW95coj10v1cwXWDELpYCcFfgzpvwUm9RcFXqhg/F03zt
8L5trkQ0j9vGMsGxOrACJcZo2GMvlY6Lxh+eEN1o0uZkZg7mYAQ87kd/GCU7odkC67V3qoAMan9/
4E6+9T9ZGYERjXzK2UqAl9/x2acOjeUPQ8Sjlw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HSzCX2rPDzjR74xLkZDw4wq5T45T35dOR85TZcI0uR8RveJ6e3Wv9t656E7yNk6ulK2MipyZW4PV
qQdhDMzhsaK78UrJ8aqkdEk9n8orDpt4scHXRvvkakLozJG+3Wivr1kSrcfci9s0N7QUzBwnurF3
x6gbVA/k1+9A48vIw1foAw5G8Z1vbi+gsg6Telm5nokPeE0kL/9yeLh81NQQYqyFcE/suGYuTGzl
DiNmNDYNJEEzUPwpbhf0EmeFQWndPmbUcYZU0I6Wc9bN8JgKhoQKvT/k3bU9EavBwjR/ooiHA7+E
iXy6nzcYZQdk9jV80EJ0zWS9x7ekw//IK2uhrg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23056)
`protect data_block
XnpLKj8omEnoJhbgAh77xyxCSWXJvND+CWuUieQ+pbgltBYO/GU34AYHGYMVmbqi0DRO1QHr49i0
2J3Oz8401+g/hC6UPB73nCOGUfCcvIOYZWqJ7cWox8EM4B1V6sRi253rjsOHDnWRFYufj0WEb/i9
4daWwrR4z6+iUA+MfGM0FazhVUjtG2DzIcyb/oJSltnhCYAaR0cO390RYZfM9zj1yKPMxzRbrGwj
8wa6hUo6y5WrhFeTqr8rgzUM6FfHfplOzp3AvDKXJtnDZsiP8RU3ZUn+Ek2JoLbxXp+8txe5wAYN
WhOAMLJOsiG/DsZ6dly06MfNIcnqzS56hpiA8pJQcD013inw+APen7OH7vJbjL01D4x6IGq03cud
Us5AvSve9yhRwGoYIqLWOw3XwDW8XXaNwvYOex8BktcDofZ7zbuYcssHOCAzoz32/ksuDqmp0iXM
sZCPYig/UtPHtg9ZzIP6uJ4a55MVcz8KSsB2UXMeZ9p+mFHkm0Lpej9YDmtfMj6GyVP5dqgGJ/KE
u+BSfabTE9Mf/P0Kf6lzJ81C0vFADIBA6omug1tG5Ukz6QWwaJ5rF94rjXB1Jk0yTdmNf4jz8M7S
4ILJkpP9ixFGPB8mPEhyLJtwLg9g2AE81Tb06ijEMM7HUIBqFlIKsEN0ITxeuKEkMoKOH4Wn9qwk
+Vu17xWrgBlVcMqRPoEqUnblBE9MZweEehzOfvqEDotZKbvcsp1wRDLiIwGvvcJwFd9Gp+8PKv0H
ZXsY6pCkr8NGHmjfzRSKK/gyaU1YY+YGRJHCv9wrc3frWqqyMhS1THnLtRBPTZA7pbKxqHlqYflX
HZ2gnHGOG2rYMHwgKn2F7S3BJ/O0+lgNY+rwoQCROjVBRZW/cLZi4o72u+wfmir+/DoPkBOjiJot
XtgxhUtm2lUxMw9eL/fiMH2b0bLN9P3hIylSaB/2pGtTa1fh1rvIzE1mQYD/4nhq4FOOrQbqiyJQ
wjVMHSrmrsiMylsaN/Dwjbj7CzkxtzY3rmjgbuiWHOGbPjR57G+eDv4fFTS6qQemGvPaoM03ZxPp
NCSB8xTBfzW+Y3DvfHdtVo3U1SLXoH1Lntr5oIpzVnC7qOKzlbX2vXehmZ8Zc7YpaCJiwnBO7uNM
xteH5kAtZZa2GkmoXYXiwYcYnE0oWyRHxZeJ3l5uRJLUt0aBaD0HNnCaZEfEpKmVsPQk79XWDBsO
oZCkraPwsXOyCsgG9HPB6E6jHjEXf1wESlwEdS1okDrCg9MCEu5j2FlqzM7CHukqoE6pWOJIWNn3
SlW2gpvUmMrgIXgRQ7wZMtc5Go9Ey1WE2Eby8UP1pDe+JVSDQiTw5aKZcGjFoKbjDStNRIm5A9RL
7twH7LpemGXMN6yHFcTNVP9GHjCms1HS3G27ps+lfls2u5vlqmfk3vs+XW0mSYxKO72iJ0jTdZHx
FGvZS8JhUI+HNmRXMz1aK+JC9dhe6unUZW8V3yiXDS/KTEtxw6hzljIa3ypFDFBGgnbHasLXmcH3
mYJc8L2bNEWEHRipVt6GRgPcoZVFX9d1IKkaAt1Jj3LvwTlz6AFEwfOU/82bWE0o0OX7XWxUiyYI
5krW138nJmyXyE19F12K/EUpIacXV7B6mD03J9FGwzlvFBPv2esyIYSFmqzDmPVRLYyT7LStRQHm
NB10lZey0P12u0F811JSZAVGxhgQNRsqggH0USsUTAh69qVgfDnOhK6Qc+0gy/WuC9E/sXuD7vZW
pYVr69Y9VGaJ8u2I2LsO7XEGyEtsBUdYtBORBKo3uC7rldzU5q4XPu5Vvax9eegeGzBgqdhw7J5D
BfOwvigOPBh8Md0F63bSGrIiO+UfvJOuizNmqA/f2Ej7sc7/8/oloRffsEKKkIXWmC8c0mXQBRzL
HMEjp+NtfDRhBbGrTXuvijwFP5e1SMBeKr/j48RdOHqnxwPbRV9ja4oa5mD79tjXjHiI6nVqDM50
RlgXZk2wRZ6Veud4CocqTElZn5vPOdTradrOV5STYE9asYq8z1+81YbygrUziTPMziG2b64JTN+g
vSRXoqzcWwEBZenjlIjNo/ojiiXSzfBPpSj78SgvG9uvCaLSmIKb6oH7W3pP4q5lrd0UtvLOifrq
acCRQKtA+9QdXmkq3rhXhtlYYNFaUnCZaPV9JtGCSNLuwnVJ0XXO8PbPCONz4NlfrRqcJqk2kJQo
YJKp0NRRfByZoo+FDLS0rTi8OQZxMEiBGHQDdHc1X4CqIL0CvFQlcAmyhiruTdQudGzoIqripurk
85GayZFjzHNa4NOmA40JQNKLSoqTAhNBloOnhGuhrJBGgP+jzLXhJs9TQb8qKo8aAVEQW+aHcbfz
FDcvQiKbCPAj33A9WIY8CrZCtdAEbJbyMMaqpwnyyhf7MysvS7VcQBbQbQPTVKQf/Oumm6u6B54a
cjXiCU0IWtmAJnEAc9SqqVY6V+89pMRGdZDzk7Att39gg3Tsv/vlI6HHlsFFGsy77rHx1gqyZILQ
R/cH8jhxoOzYIdrvffHx7o5BAKgE70SplahVucohHUFn8eKghOH6YpKlkYTDefjhAo9Ftt0qEynz
MEubo7Nc0u214KbWw0MjQmr6wpjrNdFwXLjetBFkVUu6LTsjSynxWwb6ijEoOcKit/KwTbSiLsut
Uha9I6KvSmYNsCye0Cniy/GZ6GuRtFcCNtStLxzwnXzrfl9f7Lo8PInUaQ2fmnQjEGQpyZDxcfQJ
KO/g9pS43rxv4+H0UbIODqSsQZYQOYX5O9WQcwqBKMNDzkyDvEqEM6GICO03/lQ8AN6PJaSF0/DA
Am+9MwwSmS0+qs1BhNqrBK+DDBZDQVc82VWqgk0pWiR1VxIriSbpwAxqKTuiokDsosg72UJP2etE
jUeUTELsKxU5tLaM2ISZmGDsiGGMgIAGKWWQTeZXJgRq/hBuyqxyd8+2NC3csqHDc9RdznQAdIqT
LNefiLy4Txt9J6V03pJiF+LlGg2s2DvyvRRyY4Xq7udlJA0NReAjbec2Al2QXhDSScUYq9QgmO7O
cUfXgrE4sOTxAheegwjgsp7o7CW4xDhHpsriFlgTTAVw7Uc+8iACMLtY/6LYU/AdtOvCD86kzHxI
s3p1ODYznM+bGXLfraAEdqDSY3XiB1CppMJ6VdkfGNLGD81g+hTWZ/TviBRjWXvkVOqG0cYZ2Gs1
9DoXdumuz8t2LoaKglN5QvzYkRivbd2Kk7o4KcH9DidAy3WJsf6yFGtAsz28dJg81RtW+iLTutto
jDpj3bKexvtKo8WCHb3r8SHL+5PM0INABEDc2hPnZyaw4zjUiGOeS3XTZ+sw4eQgDGsux/EoY5bE
xegoLtn8QcF3Z9MGVkmtGOqenXzwaLsXJngKN7vBXTO8NT37nncb9R5DhIkeKGA70YkifjgtknKD
NSoDpyl95+5sMOW7U0Y5/k7S4fOWuhG2dDWGgwd8Zqgkmm/kHoj7Aku5uqc5/8Z+EWz+NdKSxqJo
GaybjL+zy2KV/E0ztxH42NwC7QDgqKB7wTHUerGgye+JiZ0QvEE79OlK8N0AQQXF01R4sIWPRdwW
dwXNw/ZTeN/n3bQDgypsW9s3gBfQkhrtpxSVJUfH1uu3W0uwxBo6bJpTPxuFKlCt8OGCmVAahVnn
suXixhmqO9SpoDDkZ7tQljhsz7LNTzgUjhIk0zLz2diElSwjvNUPqzjxUAJfTrKexPrsb9gM1rLv
PLSkeL65M6za3Tv1+whxlj45HbOGJyhJDXRic0xymsni8hCCoyjvk6Jg7qg5/IKc5TfzG8qG65qV
4nqE+JBgVyt0vLYqoQ6SW1kN6mEMOAnB+VN4slRyMVT0a1HBbI0F1XqMVUoFE40UtKnO4ZI5/eyF
rejTEhqrasOfo9qGKkO2FsF6vmYKSiQotekMORrF8o3uQmyitNxmfBlDfzf12vTPNCulhxKEsZjX
AHlk7Jl96PmnbGIi3NTHauLDH9hizczhukRCZodmJAf7PSs55fU2qh/U0bobSTnSjPXGPmmJ1yLj
Sv3+luVRFTCCDfPEGOKw767oRRhvKaGcju4OQSd3bvHjnEG/vAoo+mLLTxqpfP3AY/5O5piRhsDx
JRlrRva8PjWbCP5CH/tg6H1jzXY/DlyXJGbQmEBT+bFDKScmkY4CJByoQaZC2ZyqEFQi1PL0xFHH
3z0hTjdnlERyhD4iUPcRbYLKwmXQmJqEF2KSekbVYixUl52qeWJRA4lAYwpS1drMauS1VveIZVCN
uUf4VQ1lOgEBbyy/2UZZC7B0A5JfDpHlX8o4cdLQk4cRnfUB1shq3FITuoIhyhgiKi/lun+AmwPs
FNxMnu6ctcQmS+hKcfxmgDLAPPLMc19GyRdGD1L2eUk4LmudUpP50MbpWvE38TRmAK298IFmzlXZ
nWwKsxFe8MTfBQ5y2C9ghnoy35W8gItIzG3+FLZZxNSBRljtQzxaY32HW/T0bgHkd87bcYarSBKp
rtTy7sKUpHqyT69kGyXwDgCKkc5D7mrv3yMP8KfHiwINApBCTS98v41sSyal1xxw9bkjoFLtI0/d
0WcjMSv74cTTMLIdyPUoa7RbnMwhRbdq4P2MBNnFCTKF1MejyfigptxNCUvdymcRdZ13cU62lbwq
A2FW/QWCjOk7qF8lPibIxbymKXXqMGTqiGGXSzrrnavmhmLeI7s+AZaQvsRsB5IwzMT3AUp/Ya24
hnKNnMkS8BQ/YEL/qIMCnN/8eGt6losD9YatV6j+RPa/1im+q5MhJkuvLCPBxN+6scf5thslVGpG
nwnU4RzQxCpwYCsqCGKsev+HKhjqPEJspQxj7Lbtc7Mn7D8VY+lW886eIEaOst41ygZn7BITzFmE
7/BIYJDm4/On1d1mdOUGG/+hgSLMbkS3W7BHHvMMgiSkGb6Q2JqagP6ie2V06dI7nQ8fKfc/+Bu/
BnyVvmbjwU7kGeLhxqG46hiPijuFDQYXqo8Yosq3zw5wktYhv59NXpPzAfe+Jkm5ysiOPHRbkTR9
1XbBS+YGpGHuzj2O2HI1b9NBhA8Luk7MDOAZ7B2g//3e9Ib9cweqCk6+sOQ0m8plNGA8WMZ5CYTR
jkvbv+T6wtfxzYwv1Wmd3F2SxHfjRXndBD81Xen6IGl+50bFCsM4UR4Jxl0h5y0uai4Dt9GJtOwv
sG+DE6BIjEOqzWR/sFQ7NJ8EEsTHUaInZjrY/6mepabkEh5pFTVhKTqJslM7qh3Yz/ay/hnl2Lbt
6x3HI7wTFD0jAvDuIyKcejeXP9IW1i9GVj11mW5024KadSh0IYgcrotHns2bCe8F9qrN7Hp4bAQc
QUxuGpl28dMxKN7OJKKnz+t2VmO8ebqFJfzBl1OeaIdNsIuwknum7O3i1JT3YZkexMavHBAnbYql
nhXqKkJO0n98HTF26tHCyupvyTBHfgpXcjDwLwLZEZTh4KuKdxYaqE1f7E4lu2UUYR/mDJb/RkPZ
0taJQa6acbuv5xHSt0xOeyLXPl0mvDNq6K9RaqKJXh9+iW0vW85DLLvsHsQRug7jmwAejjjmsq3E
DHNkFkNGBq1IhIs8LhLFR4jzA8dlZmqzQDmNzprQStL3GbbM2XqBjxVm82kUmRJRCEEZ7z4hE7o6
Kul6yCQU1E4dqR057ahd/B2P9E+XX7yP9IFgBYqa1VapKzUwlUIA3Tbx6Z3c0NOMY7AIRKncd9X3
qmHm5r1wDDk2+Qz5zuRndWSkRjSoD7Kftx7wS2NccE6fwJwlrI/cXX+RhKbvby0rVx3J8jfPCdWI
U6hxUVYLp7ldqPnljSHZhbso6fJ3iAYymKR2tctVHiRp7TiKpO1tChInsPPCSS+DgdoHDwgJfsEN
zrWRbcLo83xJzJbfA6C2rPv597Jdu2hCEZDBj95YIUGStsB2xrq91krPlbFmC3ib8xNMpRyGAHrM
S7YMMlwEa+RgZQfL5DH2hzjdFqcufpyUgfNBViqHy0dUtrmson1rOmB9v2pSiWEy97W/+QEIUh+V
gg8CgkXXEfJrSES/30OAqhZh0F05EvLpa3i4msgJMyUXkPzg/9BCKQaJ/+ZU3RwUlXImG2nLZWuh
Vz9UvJYr6HAa//30JhgH0wRyjhVHJXXabSaNS3/Xu6X6IBqzpt4uaI1NeGhLLAXRCR826wmIIEOF
MJWD0CZgM0HBh0BLOG6z+PeQPnN1CTy+Q/4gi9S6TkOuHil+SyWv6gfLDBXoMHQqpk7AKVLJQDGG
B011ht2HYttb+HQDSaaBmm+CMVL7tp8/41vM8qw73bTgICze+6aEUCpm4Im5vs4OVAFon2qUxSCd
ZV6wTagm8Idt/+jYtonrQTcxBghk+A5ushzb56FV5GVUOKixEd0KTxQLdvbSM4Qp+OdEY9dU1lCU
cIQwPy1TMKOL9gXp9Guq7M0Xyq2TTM7bTxk2JyE3EQbyWuSWT0HPoLG1rnHo4cQjQzDgcF5dAv+d
6tt83TWmY4khqzG9snNVUi4EmDTVC+o0UsY9NJZwLY81beF+IAAuk3gh1PVX0xEC4hogBP2IMCQo
T3rk94cY6eXLAu/LHlUgfqs3ekzrQ/bSjq/iwASaiq6G8gtQuS14nem4dvrSFcsapAjF+kJ68skA
1CktlESeRrQ4hzcUjoaGsZGuMVABiLmppGZB0EUAYLn5EzNRuojkbFXY+IeR3R4dFjjMQxpSQydF
X3qvZ3aPHwUknoXuMB/4+qjXOb3XItn2sGFuTjPG2gupR/ZJeRjBWeKbHcrvXoR/7JgXldubDie6
zXubeh9lzsgHA9ezbJiJ2uZuT+H/ihl657Dlei1ocLz3bqTFgg99kHzNyng54vq8rl4FY/HXFNhA
QO/DMo9Og6t/j4ycC7OZiUc8VfZJWykSLNsL0LPK3i7LBXf8YdpwCPDGd9VCrRUQYCWZzaZMg4Cn
j/KGN4cpJ9M11SHfon6ks8TBdq7YR0LVPwIYgv/1kddKqM748vuoVNvImkVKA7UaPpa1osEMSiYo
cVObBJR3b+q8WMLcFtt1TKC9m+rmMjEKrUQCcpMZDtzzSgGh6Lp9a8cIpu2onEMf+OTSNjhRwk98
Hr8MuQDtoxM5ySF1q/TUdKEIVL9LfFPTwMb3yezVrg9aPe6MIu6BlFIHoYVcfgORVonau/LSkjne
Y5Uzqfr7X/gvts5GnY4/6Y3ho6hsg3R9DLDwj62U6EADn455v4IPGuefPPjAKo3iQVMDs1F+2irb
bA1pkpRMEfRPNq4d8vAsk9qhEJvfJWo+xrvsjcIynK1UG3GpNEji9n6UOoLLN77pmXsvvoKNggYc
8pVJdwRQ2OjX0yWfGGS3ypg+SSTdPh2gX2lZUDIu2q9kZjnu+xR5XzRh1VAXR0CWDtR1hMpiDKiM
6FbH8ItO9IrbWLxDGBydci0EpgBSXZQzjMJGtHW5mHd0Pg3wHsSdWiXoj9M8IiuFuGBH7+wwB7+0
eYENP/+M8YCOjtlOPJAMxGEFAXMsH0xC9Uivv55jC/f2+GnX0Ol4DQ8+uBo0p3/ckez77sNhr3tJ
o3zIV8WrKVeCHZetP88kfAaQ76MYT2JdaKLYiL27LtR5hQBYj4HI+XAjOQWpE5j4eNgKnIFkgyES
OSir9nLAEnJJLEa/0+38pahL2H7uEvCyv4xgzTzQ1ysGsUITRZSYs85NA2DWCG6nSgqHw92zo912
3Ez87VXBWIXObDy/QFMVlQE4MLoxR0bCOga6ZHAjWO6CwkGQPyDnjgOdCqwuArxxqr+Rywuz1IuR
x4REaz//TmWxTyY3fAxqdcwLhHXlqWpdQ6vaBcN98pr4jZrTu+943jpcBq+xP429ZqMCiPAynFaj
Tr5hWopf003Y5NkM6tcTnXy01pLpEb2U6BCcFdRYhmkeKV1qWCV4i7d5z13nzemDGLcdE6VZWyyq
+WYXaDtxv7BVYlIsJ7hY2+6EFOljD8FGFCZK4yut+yKPZ4pVEXaf/g167lCDq13JYvHra7eh+D0V
pw16m5CsZARd0GGDnF//m7iIyk+BqYhjd2pzMLdTEr0rI6Wu3m5XUWZLMSRPifV/3y91n+3BpjDd
EqNtP0gBA2rWIh3vE4dhmbjjLodsdtuHiQWyNuNwBDl/lKsy2DlctCWh4M0IW1Lb8jo6k1pjVNIm
c+NyQO4M1bTkGyLgpLo1X7ZsPfuB3ZUDxX3Ilw1YGZedAUw4JviNLMBxWa2hnwvwQ0dsYGpQhlux
x2H7qfnvkBr3asVcJAfGifs7wN0UbR6I9MRQDWby6uNDCY5p3KemAUhUgndfbdocSEJ0K6evZPZA
19m2jn+5oLSGL/cs14zP0aqWQ3RDJC0spm0ouAzseDghIwNgHiPtSDA6xdaMgTd19Pkh+lt44Bnq
M3mXo96wbHPr/odn+yEDEzgUd1uOkLHi7e2qmP0tXGVHM/yxNFvFfm+gj7UUN1YDtg1l8dBxJRdD
FPBE2o/1dAcnEC6IGPa+4KNcAbEBJlkubFSuEaWBDeI882ujiyJ7RVR6poiwx4IwRwCrTJC1jSVt
RX4qaT1F92JsDKcuoJSvNj0AQMcOBczvC8mGoCLFhohiubi7n8ITttrGQ+7ULSxpWjtx7oEUj3ww
NtXMT0sIqBPFs1CA/YB8sKHVCGSWkKYAL3dy8hBlsPmTlaGXCsuFmA9fz4P+b/xmOTG3wzkq7/gq
8HqJVr1+uNa/Sr1/81ZpgBfC9YA6gss4nTNYzWfLCxSaJNEPuOFV3RCOyy95X6DhbBD0RmTNeX/v
EtO+/N/XEIlQ0/xGYg+kKCos0K2UZv8lXmch2Ov3fCG1azjTV7xa3OuhGV7TaAHoOJunszJWg1iy
F5aKbFYNwHoCSQAyHF0cv5Dadvj1ZphDCG56RMa64fKIZalQjp4j6p3JurLtdHUUcTb9MTV0y8N3
W5QlOzwz0WgK25cfVjUipls9J9rfIaV1Yp1zduQrmOUzlciyH/7pFvSsKsFxc/PmJZ+esx9Yy/Tz
MCWva/CsUJy3JfLYfIDn7yXC47pb0HbIX0e4Pgg90cryP9cjA5hm5WGcbun6tZd5GIcj53X+f2dO
pXY4Lf9iiw7f8bPhYmYzInetaDML+TUdgEzX/o71jQH4HyD/JjYS92j1U6dbZKWQenewQqy4P+Ll
egtogES6t/6LcpHsWrBBfanlQ8mXnlrMW2CMDsJaR9lV0wQR5v5pv3ceAHuoUa9T8riaAoI+qdit
WSkQMqu5If5a8GBm/rCogRDrvkdbtxmBzYqh8MOTIUxcYJ3fJWETruU9ZpbVbrRxZYVoGL9CuHbt
Y9Bc+tGhFGUS+tyngHCP6AcwHq7j4S25aX/BdPPq8gCsWdJMwQMsMyZbMUkEPZ1HYGUTST42Uqi9
/2gyNH1I8ppGN+NT5j8hQTV4uyhSXZE67MHFD1p9Wu0pafKMRyhYcyu4y51paQzNfDkq2xukVos5
9Eri/0q1qz9R/EzglbladEV65Cklcxhyy7BqNYjaVcOT1e6Z6P7fn5GavIVwOdUteroc91s02YCP
8U9kKWOK+52H0DfwkcsKs83cmYJQcxWyXIaeKOyHYvwbprL1wHE6dw79E7w7hfkQ2jUeKeUcMVaa
tYvrrT3eZrbFKgZ8IPy5hmQITTRBszAGGudRHH70gB/ZK5NqCeWmkM4fu181kahn4RIzL5hyinhF
TH1CTIbK7BmPL0FhhQbWo9V0tYpbClDCHes4Thj1KNJk89++jkNk5nawHEnVojDWJT+ZZ40Y9GeS
95l4T+gaMnf1J777TFt04aWoizw2oI7Ogx0N6oWndvA6CcmhTSEd4PUY4QpaN1dNRIG8HdxIXOcu
e+b/+E8rHMPhJBWQS2dKStDBbqFtUzDq8cCrvr7PzdV5brq5vhKBuSv3MybYtdpQ7PnS2zZdHw6t
qqNpLZdL2l1rT7X2szLK/ZEw7rukdqhf7qm1Of4LcaISy5ehGxpZmF5aU10ikuqM+jalkG/u6O5t
NSwZSfNz95Ww+GN0RFwvoaeXwFrZuaavU3wrwq/ct8A1jR4A1NhamuKKFCtQPltxWayysdn27oU8
OLIA6wRGeg6kUPrHQ3IVAeNvO8gFzMgyzsL0QCmdNeUY6LktJ5u1AHesUm167EMDFHKS5jxI9KS2
B01LJzzv7XrKewkiLyWdH1FCkvCJUB+ePj/24N0gP1gPS2vdv+PRMwWIOs/7gD7z8MY+63rH43s/
CZ8qfrN8VsMz+oekKxnC52MO5MCY8SHI/Y+KGD7J/DDtJgEqRxdsHASQnWzgkXWOBL5qC/So16qG
kcNGE475XeoDly6ep8Mr/IWihKRQxRA962vCijTy23DFkj1lmy5wzujHR5ZDXlTMV7A1545RdcIp
tHtbHeV3PQ3G2tLK0EhODgGBJ1jywecRXac7y4ulGkuYGzSKGW9EnmkFSG+9ibBXUQu1bL09qb53
bzstf4OWO0xv9/0HeSr2TUrzA80V7qPCc8qsug652OMBwCWYDqKa+jb4k9pqPsUAuQNIXq03fCCg
C7BDDAEschMd3cp7m7uOpTq7hevjiHWxv5q3eZQ4jMjaycYDnryI3LRlj03SjBm1hsPf4EPh5lAj
N+vApRjobaG7jOXwv5civ9gCmKrCJELcd1V7USk3X+kRowJtIZozl/I/b1zKtsP46prlOKYBSjgq
lNDznnbQ702R+Lsla6qU4rIX2g1GN281jiySCYzxJrEHkyH1wtmYuBOT3sVn6NlrGs2RMzyuQdbi
aNxrP7MVhtjREdMQZZ/gCau61Fnj8mYvlj4auvIBWmUTRduwR1V6DOH3fHSh5kD1/ndn5Zkdi9aW
s3tdc5RMVQq4pzuX8ptFj+a+H5XLp4sDsVDkzGnluNAUqAG6H68Yym36/k7ei5jW5TYcq/Gf4Vvz
/dqmi4Sz70h0PSqlMvPnRu/Bov8e593fKBUHtAxibsS/h4gE0bAoRycSZV/F0KqtpCfGx2WBD8cY
6mxASU8CtFIe6TFTFNOa88BrKlGFPmgBQl0F78LQPO5A7jfLIEaPlejoA0tUUILYKhtpQJ+5Fn3K
dqnjUddtgF0hiwQ63ukvlt9B3v+ALVr+ZJgQnmQ6dJ4rULCnqpDmX1dOk/38G8j68whxehEAVQ9o
hTAG6OPFrVgy++S7uGk3Fjb/W2wvDbfcuMmKJSka64YXyrkSuE+FJc0N+cF3rJHkxcMZGnhig1D4
haPc0E9gL0W/ZescixehfqIQDvyLq0XYmxYi6zzLdmEs7+IDodxtOVrYivae4ZQFSAGwIKtUR4jx
yAfSFO1joJT86pkbSIE27f+FcwGQVvSJzWDMVudrUH0wD7XfdSRNdL6mQSTxVKSht2UsIhRk3Q34
0b751JxjOkXh9z2yFoapdnJQrlt3knE+hoLXCFJIw1PNbX0B4c5lPDiP2jUkFlMzT4GoU530bj4c
VL2T0xPnED4Wd3oLliD866PndlO8moqb921lQrFVjdKRZ2j0S0gp478DEwkmYOT2QCauGIYLgSun
H4o81FsWrlwM/YQXq+njfSvKLN1ea7e3GM++e/BneS10wpa7S0QgM0D0eUS5NKwKWncNrP5Wo9uf
zGgaxWHqYiJ71E/waqb1QNjjtGicvuHmUaEonCnVTYfzwe7NajRzSVHEIkc7x9F+ips8dCMZyeBM
xxB6GYQWuC+vRmdoyYQ4nraf5UqWHsPFYRZF085N1TO//hP/FGpTEf1FdbS73q8LJYeQwVJocDXc
SeLamDpbheKBFqS/i+WEFcVUJ54UnsRV1ipMRXAMBBrX23D0BjTr6zAe183zzJJaMUt09yatdxLb
kD5lJOvaiBhrSJ/PbIYlMGPAPEqhczhm+UUmRy3lkXggayqlKPKXZGJf3hYuaaSxHjgFDQNtwUyW
LFJc804h+L5zt1urJ6XT8BFY0vqYmxml5IHoPNqfkhOTmo1k3aJ+XX13CVqVDMtUBVDI/MRrOX0L
CoBu45ZDAn+OoEIQAIlpNT7QmeyTRXLlfj1aNojwxsEeQf42Xe3MoRve1JV8L1fYLrp36P7QoEy1
SHV0pr4UbucbJeCjo9fcYdxL5wlTTFVsrroF2gWjxXL7vBFz9XUwzSjGVbvDN1vp1T5iy/hvF8Dy
GY5eeg0hcvqR/FQrHNJltdEtNzgDwjjyJrC5Y1pnzYrQvJVhMyVtbXsBuzmUcQwguBEE55hzoDLl
mHSdOOiSFDC26RRbxKYChyEgrVQCsGcyKLGYKrm+AeWdqzCJYMH56iJyE9wJtkjtkthtxI2q8C6L
rwTM1LMDcHalLl3zEIX38fIrl923EJTpVYwWdnVztX2vkcoFlCdWd1s3cI2xPqqmk19gIOB8rFvC
dfYZVJXTVyij3mZHPPCp1Bc8/L8vMBjqVlxlTh3JD6FE4MmtMftbC1hjqlkwJbwhdRi2hms4UDMi
wxy+jX+R5yAtR5yTSiC+brSXYMkHU5EUXd9+R6sdg9hjaG2ckeL/wjEJOueOVhGbcMV7kEDI4j2i
WDXNVZbsHwWFocOifxabhZYviVQrVXa6sKZa/M5LyjCnQDZJ6MmcR3YJKz22sQpjhunTnfO6GE9x
OVX3V3nIJz8dwtyem8Oo6vTrQIMir8TmuQrjIgJtB/6waVrbR9CXHv19+OylxZKbMFgoM6U9n6Uq
mD4VZKiXxi8UieW4M7AxNh5PEtErCVczAH0ljWlvNZOOseNNM620T+R1LXpaS935Q7g+eK/EkSJe
aP/rr1EF9csE+4QFe8twt2nvGUb9+dVuC7piGeTkJ02zH8yBNRzfv9og7b/LdYvpCqo2Omll6qvx
2S+WniY9gIP0/+ul+LlJbaQ9HCmiiK+Wi4ccMvLnKnZHpVfNAzxr8U/tNYYbdP5hHQETy6KzxhzZ
sj8Wm7ewDrGofKhdtJbKk/Wt6Yffo6PCXRp1FePoAbGMlkraR7H/huPvF3Y7u9K8MhQVNgSHwNWh
TOAFznQrJPVgoKmAU7EPIumD1ncoASCePS0VQ5KJW9IZynAj7inqGlPnodIrOVoY42P1P7eE/AtB
Iahs5uqJRfLshoQXKHDRtohPOvsUifb1vKi4YXD+xB/yzL26onF7+DYLmWieLnyc+6reK70GiB0j
wTDcq2PNpVLqozjWaoGyOTledVQj4NGzgV2/rp7KYFjZKEt+TqC4i+X75X8mKaftAhA/Bt6u+2vB
cuuhplEZVa6z+/DHvC5LqNA7wS/VDm4beUVxpcERg1yMKcDUa+QpCwXL/Ue8fUhJE/GrqCqjqWXn
yp/ikAsI/hi8bsWBhfdjTw7etM5+L49Mh5OJw3sq8/IIEAsvi/gzZZXcUP83Z3LBm9KzYsSt+vQz
5rZX287p+kWkA2B+GjbtEnoq3Za7pZQMAh1Lnt0CkSO7qsRivlZBr7hXTwAjXdE8YRrqlIxINeNa
pxeO37WOpUJO/YMCeDtI/8j256rMgIC3DJbPC2KhX1Jz7G4MZqrvlZKU1C5M0dVfCGPBCjpTNjRh
/yxlE8dIw/OCdZDhgDaHykr/7oEY5RPA2D23pMKWIVbqjA/0/Kb60qc/sdCSjqmFmvY6juYzitW1
+7Vo8MyVw/s4Z/XY9LpsLT6yd+wNrgFZ/PKOIrGr2P6t9axeBQFTMpEMCX3FKz01lr3AaNVUwjMN
8kTBfHKNaI8se0b0wnvxI6Ik9qZP6QOeGm0YY3XSLds1xV2R1hZK8uTfVK03Tjo+NICxbsBgVpLE
f7ChJHhmSQfzkx6lwI07ciF7ZNSGUw9+XKPrwqvrGWBbPwbY3KCvLDyjSU48O2zYuEWftGctrt3o
g+6GmsD2abO2Tw1fKwF04I7n2/YhlyC1C69LS8u9ZBRXqr9piZN2rrE8oy2poNqnxjmc4XKhFhDV
ua/uySJOkDqLeEeZIPC8iUZGE1dIkhuH6F9p3ai133wNDv+QW2ZV5CODeXEBQoq3wKq7UedKZqjd
eyUudNvaPihq6a4zW0C1Mf6mjUuLp8ggbvfgOCqTCa4pbZgU37EQv6rHZtxDlkKvmiYPm+ciXxHJ
oQKlYROiBdQgmPXMoXtlO1VyEn/fKMLv/Z0y0B7VdjG7UZDGrTUwCb2SJZC2CJbi3cj8FejL8Bh6
fEbw9uTlu62cRhbn6id+QOKV9Klwutxnv5PxpnKbwz6P+z6P+RMAJWzLn7Yb2cdlgGhWzFgT85sv
TgeAFYGzoYkEkIMiqQgQzdVwndmBHCGZScQ8RO9EuCIea7GfWe3hHoCUEyz6CY3TKr4adfuj69Ig
90pXuN6fFFm/+Mr+Drc1FlhK4kQ6/FM54EeOEF0rwp//jHkBJheQxyJOVt2hYi8qy/tvGERGmT/b
SCyf4LpYF9QjbgzgO5Q49aaaEpji3yy1lLxLNJN+yIpI/x/jWHoUo64A/8vOV6rJ92sNgIXwzn14
reZ1fOayOufRj+iSVP47dRKNuRITYMtRnuY4N5d7T7omMz5XuedIvb9MRuiu/xmlVV8BhpFOTcYY
rw8jg2fMVL/AJR5x3nrwnlEsxluChzskbNLyHHePNALdZhYACoof5Hc0oRGAqgb/r8Sg8GwADalm
nkcpQaq6jdY7HR4+AqtVJ558cn1+4i7UTIwFdVvM7Q9g+zLR717VBVBZ6jXs/281iOL9pqJNedi+
dJAB4gM36B1ifxdxWbi7ixp22SuDzyfViyOPFUzIQ5lMXAjNPAKVdhspMXZksYMYWjjQMDvbub0u
c7wxgVYgPpn8YNH9zPgQHrYJ3Sl2sAJjw3Pj2fOpjhR9FzKwrHJn6a4x9mtB1mczRgBAhSB4hfCC
qV5QIA2GVBVqx7RTDvO3XbA+GMMOX1FY0L9uHQAoGl0rjcRC3waNvEI9X1dKYWfU8dVMtCwc8Rh7
lAIdB3Qho7WA4Oa08sAzF1J8OEYlTajg/ymkISCQfqtuQ/TnvLex/jzHaj7yl0B40BdBRuBhTd+b
PuIl3XqkwnFFYCu4ZIwg/K1B/uV9HAMiyEIEq04Wp4Qpd3YYxGugx+fuL9zB8WRyGMC8IrtSjjC6
ql4OdsuYwtSQLc/McwaMMPDKiwWlWmHyjbWokCAoG9nH2SgESWA7ZIE1lDRI0jT0Ot90y5yeD9Ys
SGUSWNnr+e3OJiFU3pantoF20gmoYkXrr1ZCrOFU5cBQq2/qDfxk5cQe/qq4JOom/zONvr9bcrTb
VfVpX2uZrnFMEBb9xj2/ljnDgBXl++kF5gfuO8MA3eZ1aCg7l6yK51ct3ur4SX3qO45iadN+3W3r
MJBkNnWIXKVeWPa0uInkACY4zkL5IhSwPmLkvEyUXufA9Zxp8FjJBrfih4E0FrXny6WX1ePP7Xrf
xFQ6fQ+PRJUnyc3WWvEAk2SAWxex2Hdi4JtYCH0a9r4HCThAZFWQioZei6U6ZMFNpgjq+6fDbR1W
9j5TzLEI0SZWlyV/3f/lYP1Qu04+qDVPHtgjmVVLyiqmBPk/NROFP2SQqRWiKGtl2JdY7GL+ojjP
CPWuhQk6+1l29zh4NrK3GXRudW3oGM17KlktWlWbSJaDTVHHKwdvH0bNy7dBv7rXNoK9N4TQFR4e
3BuFPWmYT3G6E1uqTFGVoAQ0nsd6LrlzfFiUslGFOH66WktEOv4FPcTV2+F7zRdhtiODp2LGioyI
v+BBH9WYsX+pBhgJSqGEix3X3molM4kTSCp+hsH18WeTsPL+jX3keWEyzTvPlu5t9o2mtbcfBykk
+KpOnjNrLCCVFwBuCsfKvcBv+8gLx7tn2InZq11ImLOVgkkAyNYhGghAk5OoZfmSsPdLv52Jaj0J
NPb2ydhkx0zHGpUNPzZ41NQvoA2mepkHz/qtT83YhEieMk1RWY1F5SipPBkctcyJvaw9pLk2V4XI
JP7dxyHhmRVovsCt+1mvRrZ5A+VXtf3UXBFJC6cCbTxG1i4rXpniSi7nZAtiKmxVQdE12As3xudk
NrhbrT+kyeeeG3GUoVtJAzUVb3W1+UlJcJt3zqMscya/y0zVaTDg1qZ91+9f2lyLc0CD1hnmgQ3n
Z3NESoA9UTUT6BxER4oqSYA3NYzta8IVnA4VFf+CCadyCi5jtuK0HyiQJzIOOYuv9L/Sr+sQtAjk
PnvoRzIuSG+SXQSakiO2qNMu8horgSVzrqpuKVVk21azzQMJQtCN02fwYxsO4Y2bEXODa9Fhd+Ia
s8a0TSbwwVIJyZsp9K0aEjhg1nQYdvAYmoYXZXSfiVrk5/wIBVaCdBTd5sq+bTkSSSIws/7jKogC
90DmMTLWEXF0mTVF95e7eTw04s6UMArpe8j7fV4i8Em8DDalJHJ4Tz26E7jwntd/CUYzHh/vByZ6
2x8nnATHH7Pa7Ol1AXo8ShBaw0L0ROmwXaRFvvoMJmF1JL67EVxONvRlO29ao6XX6yfalCJN4/Zh
qfuoArKeqqQUItB0uG1WYSeM+JB6IQb5bmQhXwUt1Lk/GzfE4a5JyMwgmjVCxmZMIIKLTWUSFRzY
bu89R75npWrTturYyWXhyuV1WCTbh6zPobEshRmdI36QLBQ1H+3oodAh2V1p6FGqgjciIsm3JvRC
CCpfI5zWtPXBY0/jU1poAMQ3W7sIlCXGx4ivxrMNZ0rK5zJCip/TZ7g4S1PorUsfB8xPSTidOQ5G
gJlik2Fp0dHseI11FeLh7cRYUcSpkhPuA57O6wGXm5NR3ba35W564SSr5+B5TfKWOSlTE3//xk/M
2fEuxyKDtqppI+QSwnTMK8et9cpd+PnPWp+5O7/Vz/vJZ0Xvv0FNzV7VFKAWa+n8AwqYUamPDS0Q
2hkW+tSqKMyuMPBwMkzlkJvr7Qz0kI9aOOnAVNmDMACfSySCY2It38bP8Zg0QTmVah+8dIRYR5qW
xWycZkPPAvZKXM1eaitb9ZPgU50lNZH00U50QPc358OO+9QHOYybrJD4YCI99jYCbg9+00w6o+NL
29oRCIDkYyLMS4W3D+mHNMSxe/1Rm96ryHOPY5gQOfClyRhgqCsetkYL2tQiFcB5HzOaJ6IW0zwS
eXj9xsdP/3No7au+BMRjR8VJgDGEnoPXbTFU4piDIc/0FLb79dYvhLtjiVv5Y6iIfMqt01SxUk5d
yRhQf41JxoRbLvRSKsyzAb4Gb3m53kCcFQYvb0jN2l0pcPec2YJEFbDC4cq/Mn7O6n4Gfm9nzQTf
iEMQIW4cd2g2d0L7zDiVnWhfEIee5PShVQqwkooxDQlmQ7LbTeuaMhD66FA/QDmrI20LzcHCrklS
kqseMYUH5hLF0FIm5fJqQYy22lz0XJv07DXapfmTsOsxNcPvU0BEGBdpARpyY5VukdCT4ZMKIm2b
VxbyWLJMnQ/HerWEbR9yDfsPDaduBbEp7J1S3KHbwXmtGOvZ1OIw1zexPkLKULvPaiO5boWqQFZc
xjRfwkW7U5+0BsTxI97v6qhw4DuYlT16eyOH/xkm8NIVZB0tb1iA9pNR2z0fV+J9J1TigeL/+1Po
xjQBL5g1E7WHmrq2Lyg3ZWozKCkOPXKKsaw2X7zA0sdnSFnBgk18fQkl/5yC1HfLKivN2dG1hVgT
2A0R6BVs+Gir2lvAJx3PnMwIXQ/IXZV6r2cDX1sMItp6MgULmByzZMkBd4Tp/xjP+zkfwc6PKDLg
0bn1c0v9SeI5qVl2ChRDH9DjgvyxhUJ+1Jj60Ocujgyb9fJ/PSpV0xHNSL/uJ7Hpm/I175/HXYFy
fHJV7QPX1L1008UwFBfCm98o9RQXsPVHUpELq+gcVScgGnF5VKaWw7zQWlUmzZQ7uNwlaWteZAll
Hek2yIOAhpbl2BxbwzMb1Tq8LstAH5yB2+UNrSAJprUhgcaAZrLTpF5eWxvtg5pyh9MTtuZDyyyM
8U1MqG4DEgOVcXS5ITf285u8m+MAW1vTCF8lcU3ekwuqbitrHQK4P0tLBrLJvjY+TySGvVwOY6hR
3Y+0D0wH0ELftu0wA+pUkcJFN/Vu48EVx2MGblbpvECseX50N7KcVeKcR//shzqAfdnsQaLszUQ0
DtRloJt0yLPeiCPMGQbFAWS4O7Pa6ulPvhvp7H1W5tkPh0i9U/1JP62r+KnGDtjjMEsidWe0y0qU
wbhgsuooB7ykr+rds3p6SUY46X+ye7pNygkdbQ47JS7S/PdVzzz6K1whiV0h5W0XZC7g16eHAxWX
aBVZF3gZnwRdxfH7/JyAwI9pMroooGRDlcE+8qy5pDbbE2sIcaAsQS+tR334HDtTFW5n76Q2FHP7
vdq77dvhbicN0gVaYFUfe8tnXYXgCBxm0NTexyFBf6aW4ysOCjUx8yVKq8Bj8DlkzsALIhfWAsIn
Pid215bmHfZCfUTVtzfsPT2NOkZFl2oF9MWa2s1oomTzu4Xxxy+XTA2gt9JJzmdYU+CYpJthWj53
eoXVVnVC4NLgTTCciYzOTn1KPhEfhlLcJ/1n4xuk08Xuo41DXs4RlMGhc6WFJxR3ck76ItZSnnEE
Z2Fq3CjVjBCMOqoKv0n8CamuySqLcgo+M1UXvq8pjdz5Q1T3/Olf/rb806/ziltiaxE/0iFxlY3F
KZm59BXqxsCPztgIc+0WZB4RvJmJqKoRfv5K5omV+lRFQvI/R5k3xJZO4gwjFsAqazmEdFRiu75S
I5gDJrhLSwx1JjS29YgaBjuhML85J8IfFVtvLIY5nf11pV2S+KwdMXDwMWiFdwgrZcYvCiehgFsI
8EssgnAbJ/zIzyWshz0yOu1s6T3vRmeK+brDKLjIM85zgyMoBCTmJBukwdlhSi/K9guTIT0foYsy
S9AXCKo7/p5mFELNchQzmrQOuyo2ME6j7K8c6DVY19Y01Ii1Akk+tdh6qj7gWKz2ytV8b0Z8McKB
QHg9eG9v6qET2OxMWuIyh2/p1fPbIKSgbGCJLRD2esaE9qj038F/esmOwwQcDA31J276TyWCqgzk
pyUBu6Ekvff7BpTVU6Wln+yAut0XoC4p68Idv5OERJ3C2dmEouneVsH9O++cSc5QGSYGDgRa1s83
EAcrnfocVZqhgQFfj1ElSzxKiEnWC3x+5O/rvuEQACrSWVQP0M+nWFzJWeo4ef/F+f2GkdQRcDOV
9ijYWHEIXopztMSWlhJJi7r4iPsEI1vbc+pf88gYpKmwzezQ6ZnqQOx0RasFSSC1uNlCvGooEk+W
RoZ6ZMl1tUpSrzD1HEDmbZWqY1zkYmg1F4/5DEXGM8wqf+X3InA7xRvR43zZZ0tSwghw1d04bd6R
O60pEXKP7OQC47II/EgtsFtfx01SvX7kuJm4U0bADwwnEKo9jP3HwTOTb/uwNaO1AzFJ7gWMwp3m
ar/FErxiotskJfCmx0UnfPEujRShcGQs7t99W72pMpR9GA4UaGU7vDsetdqauk/iAM7VkP+gshnc
z7i0XC7bJZVGx0jXAxbq37encqtt/pvTNhCs1A62ofNTk1s6BZBsi1EOD55vTwXavW9/1LHmgMxw
phsQYJAoV8CrmgJwbwjTczepdcrvX7/nrY5Cmq1X6TDcqT5YUA0Bo/jWn1GHswo8HqjfWhzz5Q+p
D+doG4y0pB/GDrhlGM0z0Bw9YinGtoecVUjqhdH5O2ETiARn57T6tZm97ugckayy+Xdzv/da9ePx
K8i88Oalo84UmrlhKtscQTHF0p+dWl31OjGeI/jaf+59x2UorS29ORaovjL7ffi7OLR+R+IKXG91
A4Njy2CFZosVBbL8hkqDZqbZz3KskMYXxb8Vlr3mVhDrL1d8lSR1C/XfKlekiE7feOmQyrfSKk1/
Iqo8c7tltfFMjHeend8+SvhvLxBfbqWIKN4ehkdbjI/OTFYaNTx9w8mzUxl68jLsj9S1V12DXRIb
h+wgDAk0LCClcGjU1rlIhgTOQLZOsWy9xixrh+pooG2cWHfaft/MFe/P7KwUwhJq47ydAc2QFEcv
om7yluqdz+lH/jsvL9EoU5kmTONphUygo/ZjJ5xPCYIag+/M3168lj/8w5y84pZ3Oxmn4FPF1TTj
1/33NGQhRTiKigVqs8ANWXDGFywXrAA1zOxnVmQlLJsJi8i5UL2yHJs+JjSxkT8h4ewh4SVHXGEe
PbBWYnXhPeOnpAmc8u6HAkm8Q5YsaoVptYVVldtzHfGA+sNyjpXRt8xtJjx9nwdnabH0vXwRezth
rp2dp8Jrb+W+jjhZIPp7JhUuifmnCXGxTcdhqd//7Tp9aBuDsJVXrzEQ62S+r/CAlLxqYYqyEHXl
As9lT6Ks8kO/2mu75fCZipdBxV40du6GKTkm8oEw2/flTWY9Vzet7ZDgjlFswVfhydbyqbmQgjOq
dkfXDlvHS3IZJy16BN+uNokaGz5cJbzQbpgG58Z/QNw7sXRXweTMqtLXIG71fKUhpHqyhPEDdRNz
bSWJ+4tSmo/VxYBkRLBhxdZOYcRWTQq9RD8d7Yl0K1DaJRdGisEWo9DSa9AnX+ooRYegnWThr1ec
Y8mH1ZZT0Lk6VkqMSK7vQuy46+K+4111ezureQhklDlfBqUuaynbuz8PNC5D/dhync4f2KXyFqEV
my617lX+1WQ8MvlpzGuGa+kmCO+XXPEf+hzBT/lFp1gao9l9nK1Nd2/pLegRYFYJwDEQvmPnhOHp
Vq7tnHOId+642iXaH0EzFoZOcG/MsHFMyDS2qKKihm/jVjHNEZ1AQnnTHCscbsJvjbgDA3Omc6XR
s+iGJBAVbSxVY/jD8oPq1kGABTMd9UibPquoZYMowuv2YDryqbKB9hVoG36ADaFTk1odrb8vVlaa
fRa3zyKXTYMhMHOmlNE49XNONsZB6JDEu3He3VGUUFTLUlLXLxdeoo6Ui3nyaAysugK5TjSk7XH/
n0umIt0NF/WYkmrAVs2opXQXawCSa0BWcIfVXGwfnaSdQxfVAYwlavgJLlHgWoRiF4QmSPWsKKL/
D8uOKVkTYhDZKnOzC/Vrudk6YwCHjmPyPvKcI0zWuKgq7EbpxtPJP75E7SkQFSsm8pfMLdC9iLJp
76QBxdj0M3d/Zn+8u+rffyEoxu4xF6mb0kVuowLCvFvRwSbPcHp9rE1jWuBBubUX54+1GEIlahWf
//M6TPP7BV8l0onE8uSYUXwaeZ5cw11Q/Onko2uzhtyBJXdgk8Sngv8Jv1eGSr1fcpu7MIwuHw+e
YKFmvxGbb2+Mv7NeEIjKTkkwv3Rf2qTGeBlwd3zonjQeDqtSDdN/SERI13t/g9luD5MsPUGFGqI6
qJC64cOHi54h1uhBF3/XSy8tDoFWrSakp0dDfvQQztIvb0lbeqn2XAEZLmyh/6WlcVO/cpVxiyUj
6uw8Xhz5Mfo6rAPtaym0j+LB33c0f8Y6A01fKjMuvDHNECaohzQjGDtk6m1ZthavagK210jbqow5
Gd2tIbuDUoU7nUVlbZ9mBUc9so9oFlC+jT8M8LCltMyFnrr6ucG2l9uKK/mzXdDBdDzl9lXRJeEl
PRC4P+sNzG8hmQsAqZWqiZdIMFsH0BDZNUG/4yd05VIXi8LymjXvovAxR/jS0/SpM4I0/6xT57xQ
IPzHQSlH0NlA79h/yzB/vldVGgiZMxj0b40TrG5TycwW7XR69x42/I0Cd89yues7LPCvBgmx9OjJ
xf8yO85Um2Bk5Tlia+aWSD5zDTmLbs2ryrWne6mnFa1yW4GE5+UFKBNEnHovpjban/sPv+7R4BV0
ekDI7F21RZHdRFa+g22O2GBVoQsj6vu4HsJemh+NEvveFDgWtP67dZNX2sKoOcV3VUPipoCyhTCK
H+4/gOfaO6BWTX4EvKjxkUm1Qe/rPd7+JPK3Kr3En/BZ7SsaWZzTRl3YLvy2umGnT1Z+xmmmZOac
/E5XvxMcc3qVpwshmDyUEalHYw3RhVHcb803sy1PvVpkEbgLue2fhj/OhAkKY2SkB7Hc7sh1uFcn
KJCFHE9qVMv1Ke4QVqwc5uhP6gIvmQm9ckkwApO8F84EIDp+sJnu/wyJTjj/ZHYAevbmG5ThCpZJ
qylEoBLXTcmGzAD6Zc/obxe3stfljEwTY7GHDrzhjyhUalijFwBifATojdudfZqP5N2RvoyJlgTR
LDiaK8dbH4yWko25MBX2SDaTKdAgfz3swtYn+FILKXSpuCCMHk2U4CnlNLZMptz+Ni6OrMV9kqYF
9odEA6+p6tySup4Pkvcn9zqurhppmry268upehnLdLnpVSWyQahAaIOKoZUlQhD6N2VbTy169oJa
g/6FxXNMhNGZfZuiatpuJZoY8NBzk80GLXfbvp6GBpeUfF5f7fZ2HWHzWKgAekZa/jiDZbk18P6a
/glME3Et+1Cyisn/DqlF/qzbzGonxNCmHIoXQ/Ps4UQvdM2u/3FVdU92nwqUjAMg02XTuYrEHA5Q
oZlPa6wazCRbAjJeoCTI/3/yB2NovTS+XTXhTetQrE+Cw8WcEFJRWh+qe0wiDGKEn34FbNZev8n+
vLcqWWURoBxrFYAnXXL0Wn9kqPv88+5butD1FKpbanFSeyTtaljjnqk7yRNrhopVtTWjxsNimR2q
tqQQ7hX7/AW13G6pcXiS6R/rG40vQQhmYSGVoZTKWqhd9+pMA+n7Ap+5RuPc4thA2W7IJtYZdzDF
t0uc5GPCYvQJHXjFR/tddQf6cpGoEkNKf5XmfEIGa3eP/dBFsF2g1Y+f7/x4pcyTDzKuqZSzMWbd
WqUV4yTXr9Ec7+Ydepy2yKV9ZUd53ivrZvmSaLZu2FVRyj2YLoHh9sf2gSmqIky4gTgkW1a9q9Pe
Ie8hZKaGCuVSkvFN94sthv48/7KBv9+2/OmFHRyfgDUWW89tmNtn9L661Hocd1rN2QFex+NCAfFb
OIqlHDz5ouJNdc+sCxYXlVD3G2cok3uuRwe4QqMGP7bzMts0PAXB6q+el1tMp6DBxSCVU8+Xx0ed
tm6iUuBc38JNY1QeKmCQJWaQj0Wg9BXeFN4Wm1mXwxJ6+clY2fY2EP45Stt2UnlMaYjod5Zu2wUF
fgZVY9VXjmi2uAjjytowfyTM76PRmtM4iBMlHtrj1BirDKGbJn6dZZptZF0Q/Qqb9jidGfU9SNPv
vk7MPGqniTZJRPW653hvghT7BNivC4KDMvksnAM5yGPCYA0Jd+/jD6g/eTa0tzMA+sCx92Lk7ND5
pHyMdsoPmkXi01hiV+RyiAnvrcEHbJNi+VAoEGB2GyYkyQ5RtVWuctScyyuOxoQsFaFgN4GOWe5e
nt4f9QbcWQjAv3rpz3Hv6bWcGatLV11bIYT6Kn9N3B940cK+TyxdCJRU2v/Vlia2Tqz3mBirSa9U
kbrRHUUTnLodLUHnH0CsK8KbCA9AH4q3/Izm0UI3tgyKe7YC3ScV8gWwZDtB954xz24aVzgX3KG+
uojTrnim37zCuOUlq1Dl8/TBulGHIfRCTU9r7yetnNS89WvGV8GPMAlTTW9MYDNLOjpfskaGGN5r
UrbQRhFHMvoxLGEOzQHtdy8Qrx5OcGYefBA70BjTR14vzvlgzlsiWvME7BD0R4gdIVbvBJjjcSHl
UCf+cGfI1e23PNBbZNWYe/vTfsH6K6N7Wa3a9Ye7AWbb5DnR4crAAA1rsGt4KE4F6gDGJpy0fZ1s
/ekj14v+abREP5d/l6ixXgkL0/jbInOlSCwRNEykzN8hscykS1VN8Nt+PmfBTaQe1sclzbBRWQiZ
0oU5T29J88q9jX9HyJw0YwNRu0RTL6Jv0kPvTeJhbweCOr0R3rTJ9dkOcXo/jpejX2J+W2UPh9cZ
Gneo7d1Pw8Y/haP+9KXoihHivdaKimhSfzZPGAOiarBKqrb1AjR+hcDT8KUKEN9jHUMCPnPxW4jv
S2ADkgCzyRTEsBwJDXPVlCE5dDwY5BpbcXBcCmerWZysXB+ZN/aOiSJGwWjLFLXxK2gjg5MOIqfH
r/vl/ej5dLI7G7ebAdUEVALUaQNCurhH3M3zD9msBRH1zMuRvIK3621ACKyVsW/laBnYFT/BfSk8
4vsQYPfcuWLIJMMRjWa7PpiLXLsB0C9ZOEukvj9px/D9pBzFCbDIj2ey8qIPg9sWQ3ZwdyEFivSb
PaoxI+4fr1xDyeT5wb1k8KO/sVClQay4zfljQFty6LfjH71sBEr87wuv9jbJ5+BIJ/0/05QTPiex
AzqTR1a7XOwTkoseBkqnnY4fEDHIwAvWeRnY/SqNXuevzKBEYtySRw3rbksmQhG+o9aMsPFS/BPq
QMo32psBnkvonXDLvoT8xRv+9wDMRbOXOHzHraNvt1CtXRDCivPIoiG6SeUsvjlferZyPg6tfbuZ
hVeeoYnscxEpC3r3+DpanEBlbHhwpy5nrGVg4xKq8P93HXaKfRMC0/gQg9dYKwsFH133eBk8T3rG
7glC+3/T1WjdJKVMxIkgeuzQB5nrBR1umuqamm5tZzpIvy6UZ0V9vgnTPmmIRGoMmlSnwio8vcNT
Y9CZ0uPoxXnZOUsvQb74V9Ksr5OcG8ccCsQNNr3sEiV27HhG4bY9sl/RZUeTjzRCsCDxdqb1haiq
XQb5BAptl0LgGm9RJByWpKD+0TyQccjETtCqDNVVcnRjRSUyROv82K4AA3iFzjyQWgDIUpV/DvHl
NAuLgn+aTdg/PIgiG4+FSBPMUFfPeiNRNSEKo/odWGiqpUjna94IbejbgxXvFwtr5mfRtBCv6FfN
VoCHFw34loBzCLsAsUSQFMwM51z6mVZsUTuzLIRXoATCW/zD7870fBSNQFYgCowjLzKXfrB1c0xq
BRG/FSYAG3h4p9435johConE5Rpu6E27LFncpNVZVaMGDD0v3X+Bc4LZeN3zt0UNUqiadG77Zs/0
qkfEbrALWpaDcRXppmcL5kAqx76X3m0HZy8XlJQlQnyWI2E1sfHMagmW3HbAqWPq07QtGkv4yutX
rQOd/YcsWrns0R9Xmvk4sV/vFnRv6nmMswwygWC4AMwRF49J4atS6TBgmBuoKBXaGmLtqgWbzs64
32nUSXN29FQ2EkDs7VI2YP2ZmNDkEuGj78qIYJQfLiEW/FFAlMN9fBbF51G7Cr/g77liW1ZvAwlc
dZuXPOU8X4Z9iaHH+sajo45HHEOho26gGf7AzXy7sihLqdlFlCRsTYbcI5XHx1AESqp5qJKKjcpz
V80CHBvsPG3CkmQuzAPxbaoaCDPpPoFvUedsC7wBH/qqVp4p5bgYEe00FNLLeZvmHhNraXRBsyZR
IqOxPYnCXlGdfNb4fxQOJRep4aJV+z0tdz3aPe5G1pZ8tI5pc9vP/OXJ9/ebFz/NO7FKM4tJfgNG
XxMMG8VaSQGHc55L7crEeWdsscsGERkmdEGt13UaZ6H36S0wlZo+Yudn9egUDuAze+qndwEQHnbl
S6yygC3rW2TcETkhmW7VatXtkIZG9Ji+H3aJuOTEawdRtP76d5dzzwssbv3yS+b2PkgafP7r1sE6
HJ+zQT/M1GVAhSHy91qtJRVufhEzfRVcugNQrgAn8slSfkWCyKgL7n9UOrR02VlICPFLMFZHT8O+
eJ8m2a3ZjS1YscJ5bSo2b6llx80bOs4IKmnE+mgt0YB/BdXAHWaUxoT+gqv/la/inMOne8JWmOcj
vzzYYJUz5D5t4rIGax3UNA9/ujQJrgXpqj1ztn1GmEQbVin6F41n/M5OtXY9Q7OFyMEdQ1tFqPv0
d3z9TMsLeKn6/4zJMdQ61JK+zYvyZOouF+FHZLmi01sSrhDUhXcB88+YitQcTBU7mfOmRmQCvEBg
PnjaJ/fb84HP57rTfPXY+CFGz6cEg8xHBrqAOA5fr7iIt5lXb8hcLMcWVoebXq9/OIlCoUux4IU8
gjVQv6n0tlnZ57HjoEnzhS1NnyFa6sWvT57ZPgLTLmxvEBN0UCCeZgLR7q2dP/NkLpiuR6txJFKm
xrhrg0HoV7mS2M1g0QCpWbN72WvlVjPTCEbi5FGlUlMwoQzvFo7QzgCgCesG3fEJ/m9XvHbOg7IJ
NYK6UE0BPOvfPXY4CywvhorZSSys1nKRiRpYZuQLMLQ3+HhzGzXs+rQehQQiV0xddfnRsDxIhEag
JFQWEyyPn4Drif78FEYURYs4j6pkCXBzbaq6IZUfV4gXHTqXGkl/nXDbnAYJ0qxxmYanI2XixmK4
bAekKrt+TwW5ATZtMgmZ3A+07pFNgEa6nbXISFN4YSS6ZwzyAy5EBJ/L9YZfZhaUWk+lG27iHEPm
59eEgcu69OCIl/aZadF356zlhMZRhW2x2jKyVWeQ2C5Yt2dZ/JSD5vgiGMgutDFpY5DvjUcHwjvA
jeK/bnFkXLLxOvOuXx4dkWEpP0/BqCoMpTKqkh6lsOHVh49PiL3bahzD1A7+yWWHgJRc3FLAhpQB
jVfTkq7dttUUDhQh+z47vq4QBmdTd2Bn6a7SbX0GZ6jrFqXhOXfPj3M64ujy+hhYtuKl2DbGaG2W
fy8mEo+s7i6IzxzsmKZdcNS34Y6GTJbCWyhuOZAMNBVOaN9uhbyd5dCBsPOmGVIZFQyOKDw0d5af
BQktBAeHeJlQo9oUTe39isaWXEpoXrJ/zzfI+tzbGKdFFJ/iT9zbbDeIp+NISXRblrjtmfWepA3N
80DYCNQAvtO6ewsfXgU/H2TsJ+eSCWZSkzJbwufPhLfZGO36S3fkNHz8wx2+KiqRcjlkIPo6Sn72
0FKAnk7xXTOaIOO7VNZo+OQSXtklpHi2UWdqG7VWcE++9w/i6nGJ6jsqj8lYme0c+gkIkcpe+nGQ
oM6QTToFlLx+JC+GtRaVJYvOxCthhmFSuP4+voWiqCntqqB9NQsgYlP98WqZ6VUxdEVV32U8SDc5
nPAKzBOce1LxJjT5Yvb9KDhLo/QAw5l9CnJSiB7a8qNvbdK90ILkEq/sx/vw068uTrZAL+IL3yVR
PsmcLs/4LzLpbzedneoxKwcEf6yQDgXJiAwkY+TOSEPxcJVcBYACLyAqtHYNxuaZtoBVmx87ukAW
0lftXYOYIaHrus8BcHw2Yhv0/Y/8F/hjj2+1VS2kuGNPVlmHbxW7bAINc2BOuXcbOp83wkyqWCUM
1QRtD+dznB4g0RLDYqBYCu9E0lWh/u/zLdLF+qNOeR8YOE6SUfgPbrp6HWTmpYt2LyD/UVLSX6iA
xC2hBjVLQ9CAqWQSarzbWsGzUsYxHZ02wgGXTbtecVrCE5Mxp6hGWkvfhJrbsrxDURofZzeNUqNT
QtK+Ut5jngR/sHijok8eIS+HuXkNfOZMeYgV6I9/12wN8PalYYMEyib4Y8APXdozIBUpaU7kxwnY
599hpMItS0StdMD6kXE29I/XEtXzaKnsiqoyB+Htp9x5o+MXAG7KMSIwm/f86qT4Ihe3aacuoTL6
ybkYD7Alb/52plPnaFwl2NxYTz05hWRc94N6Uhe6Fk1ysH4hB2eENaQM9jjezpIYdh+JNugQ88Qe
Ab59eGljdU1oQCFL+2VViJyiQ15WPEWTJmVZ9F3cKn2MWgXnu+EIKCu+eG8rQ1U6AJ+nT3EXRh6C
T0w2BFMzRmzGGfs9wyKkFmvLZF2oDMVlDuIRXVoZ+Rge6Zj0fguaK6VaqU5T8YBHG5j+X3I3Fj8E
QDF0lDI7DzP/myE2EFMkA/HlpsRhgM97udVfk+QRw83mnN1r+veCCu4bXNBbN7vf0hAmEW3XuZsq
yg8TZVntyTeK5oc7KP7/EFi66vBLinuXCbuaHyJaMwTHWP+IJRaf28xuoQ2Zcw9SxscmvxpWU3Sn
rS9AfLyPTHkvF5ahuaCFFO+hDDCUwmBZooSJqvIeK4dZfmSDeaSyLBJ47qT0YBbSWLUVkxwJXK3O
V7U5SE0qEMC3QPDp8+dY/Y0F4la6kvs7eaUfnllHDH1m3yML1NJzEbv7Z0R942AnChJZOXqdQmfN
BdNLBu9/J3uy7csyzPAXyYLpYxdJfQIgb7eyJ7WuhUuENfowKHHTFKxx3NxpZxT/nFB6nwR3o/xc
a1oeUZMgfpTQNeF9/tegxyOkq4/Vk7P73tg64AZplSF47feQDsDLbGO2MLFuoXbpesdaZrprJRWQ
uBR/If7lghVLrBVo7sb91T4fdAllrMU9utm/fYoi7ETY5ELeMjyzobeVfkxvAwzP7bwFMq8JiEm4
KWmadQFKZx1mxT0ANYth1gStX/tIkW/YjQmtK/AGSrRCG5dA6idGU0R7CqGnb2XuGh77mLPwhPnk
JUInwG6ZpAtw7iARiLPy2zWOB86NYrl7K4FRXXIFASBcm90S+67hQ7YwoOFGMXlra6lQmlCioSZh
YhdKBVoA2gaj4VbnMWHxKFGe79IaGUzinVZW0Ao7mGjRi047VBPfq7spjjsCVFRfVk4SEFIftupO
LqbtG/Nae2EalM7gzXR8ZnFW6+sxIwTWVzi+sDcuiVvICdnCV1ktGrYuBEsAsmLjLtH8OTOl+3Xc
reTLg3dSBDUkgWLAfc01xUNSPPrGVGMEgVykr6QSDJ9dl7CaOx2RtBEojmhapfcXDkaPEfzoSDwX
ZNX3a6hD/j0eq4sEqgO5mOCEtB/rOmFXeVEvFqsQl9Dn+OQc8EbnerY8LYje2ukZgFh5z1ENqCjX
4zSig20A/ULmp+pVg60WVRg7zHd5F6uhXQ66F+Ag7keNxwqJ2ZxfzXmm9F7bUeIgNHkDFZNJYPyF
eoV8DFOL4w9+VXx7s8OuQbC4f1mja4/smMu/FmbfH+WC5XF4ew4yQQfS7OW1/9r5aaIPdlliEIez
amqvHCaHpPa9JWyjhGJ2f/y7inCGTDf7JdoE+dXZQpXYTuIC06f/1ifPjs2I6rl4v1NzS19d2kFX
ps1AlLfLkXz1vFuFOA6farN9mkVA4gKKbeqsVly80ZtIQH5bq546iNEBt2Ya4EJWSTNqyuL4fkZR
OjjBOXnTTXFmAY0ClbN0pgOsFyY1btvEpWAzG3+ssGsoshj9AlXd0eix1TAEYl5+1FlwCroI/6F+
4w/GZgOzMUYkGwNcNIrO0pfw42SENvEE8/5sOzpDV4LgdQwLe0MYptZIMM0fvA+uiUK/iTn70Cnt
XGprWUT2Q1mHABHl9CIpfyDYATrWMJAbtm2tp6WlE4xeS/95h2Kjp2yPyC4xjxiGGULlO7jeH1Nz
Ze1TwBg4ulqqSSzrKkZU2AP83c0esKAA0UiGLL7/QdwTg3qe5h/Hy+Q+3vfpi4entNbF8DJbqvr1
PvIPkTs7yCy4u/DjXxazAQ/sS3uiqeFU3GIXgSJVEx82EsnOqBmYMnKvaawxTX0Du9BFYIsMCWhH
1eDvN1FjbPjw2nkjWsFbq1zbOJAdVg4dXheaJvRLW0ZTCs2L/gD9vBRmOe0S7/symZfdinz0tloH
OrwyTNx2n6BVk0BABMDhoJRqtjWn0iBTPVibpu++kYwIKLavd9whhn7GZ2mTnc7r8ji9+Ig2i4Z+
a6GM+B2FFyGwg83bU8ups6Do0y8jKwxTNR4CvOo8yAKLpI9LpVMr3JdS/vk9G/cMIuv1ab6pFb5C
pLtk+XNAQFoBixlvM8TOf0ZuUAuXkgmBkaQeDrnBmpsxE4km150svGrtsOt+RGpDy1O5LqAq7+Mi
zFp+/Fwd6WvxyYRrQMyNcwAqyh8llHEok9lhdQAsl6DSuvCPd2+ymQUQqLTO6XeZtamG3vP9xFbb
rMcVhqu0mHHIPckW4lZEDM3YsYuAcVwFGfdEyrz2ijhsdD/QWUgbRLQ4uOYElkEEMcJxLCXt59CT
5BxSRmOMdAL3GsxwWEFhE0Oo2YT5FA+FUjBhPvynLuu07bMHgnUB4oYPutsLx965rg0LGA57Y+yD
zrmDyutKrAp2iXvLi0oSeMlYkgfUmcVcihKx882YJmo7RCrdr6F1mu8u0eKqoCgCP/2a07tFcE3w
jp2fhDswiFOZanHZIh6mtwwGalL/y08XjLMJ89+r4Rhmednx3bvAxh2ucHrnwivUObAK/r+mAqmm
5AwIh3LzL9yOVRcpv9gvQvzdksomWiMmylRUWCMFDFwftsi4YLa0fPKygJxz5TRCx5DndH84TRD1
ij2miAiLOVAJTHCTbMvqGdRcSS5oFRr0U7qK5Jpnig2vLx4shycq4L5wZjT0jun/lmWPvn6+2q8V
J9dC4RL4uTVKGPWoalQTgyXJxG/I3oOS/UbynMyuioPnzgELRrQh8UxwWgqPICKFZFFuIYuu+AUu
6NtipfUMx2VSHixR5Lr+W59y25hJ41o+PrXh1HbWr2OUD+ZvY53TnMU9HKezcrO3PioLSvnrL6IO
ccASgEJ1gdCFhB7p4d+5xOUwH5H3fBv/p2M7KiIw4vEpg42u96McRD1BXupeBY21eTLIHmp6xLIc
PAxSLAGBKGP0S/IsqGjwwSXZcfHyzzjKZGSjfYFshSRdd+dnOY2p4ltcUgkcFlMCPGl4+2ENgb4Z
KD2EcZ47Jo4cHW6Tnq+6UXGh8/6/MKJaIK1PjXiUH/VK3UGKhWKqU6J88ZS98+6hkBJJgecGsgyh
5sUl7v8qvd9t/nSNriAcCkBibkZ46zGSY7TLCDlrdBI2ybBmKxYrmmbdFEOFt6LJUtVPNikBEAoP
wDKVohN3dfZOkNjSyqzxLOJpjoaTEKDOx28y/YutHshq+Bj/9bPa65pLDFClO39BFJ9PZkRkSBIQ
6zia/m9JNPI7UuMpRRme19oGBNLjg65MS1zGIucYWTDcQOCLcXZ5a1q0lCEdWBuU+c053qKOs2f1
ZEFhv6I0feW2JJCOiyXw2dIaNZaxzn1DVHci8ZkcA7fFNiwOYFbjt0p0/B2zWTNUGSzXP9/vvz1D
kdLazp+ilMuy9oosVddtdPP+bkyxMzZNBdf/mOjSnmFE3PTP+JhC/GvsB0rsYhBkWEt2KE330tnA
pFmr4PheRMeYF6r2/VdvgWFEwWNsr7AEjmORYw==
`protect end_protected
