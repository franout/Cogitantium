`define NVDLA_FEATURE_DATA_TYPE_INT8
`define NVDLA_BPE 8
`define NVDLA_WEIGHT_DATA_TYPE_INT8
`define NVDLA_SDP_LUT_ENABLE
`define NVDLA_SDP_BS_ENABLE
`define NVDLA_MAC_ATOMIC_C_SIZE 8
`define NVDLA_MAC_ATOMIC_K_SIZE 8
`define NVDLA_MEMORY_ATOMIC_SIZE 8
`define NVDLA_CBUF_BANK_NUMBER 32
`define NVDLA_CBUF_BANK_WIDTH 8
`define NVDLA_CBUF_BANK_DEPTH 512
`define NVDLA_SDP_BS_THROUGHPUT 1
`define NVDLA_SDP_BN_THROUGHPUT 0
`define NVDLA_SDP_EW_THROUGHPUT 0
`define NVDLA_SDP_EW_THROUGHPUT_LOG2 0
`define NVDLA_SDP_MAX_THROUGHPUT 1
`define NVDLA_SDP2PDP_WIDTH 8
`define NVDLA_PDP_THROUGHPUT 1
`define NVDLA_CDP_THROUGHPUT 1
`define NVDLA_PRIMARY_MEMIF_LATENCY 64
`define NVDLA_PRIMARY_MEMIF_MAX_BURST_LENGTH 1
`define NVDLA_PRIMARY_MEMIF_WIDTH 32
`define NVDLA_MEM_ADDRESS_WIDTH 32
`define NVDLA_MEMIF_WIDTH 64
`define NVDLA_DMA_RD_SIZE 15
`define NVDLA_DMA_WR_SIZE 13
`define NVDLA_DMA_MASK_BIT 1
`define NVDLA_DMA_RD_RSP 65
`define NVDLA_DMA_WR_REQ 66
`define NVDLA_DMA_WR_CMD 46
`define NVDLA_DMA_RD_REQ 47
`define NVDLA_MEMORY_ATOMIC_LOG2 3
`define NVDLA_PRIMARY_MEMIF_WIDTH_LOG2 2
`define NVDLA_MEMORY_ATOMIC_WIDTH 64
`define NVDLA_MCIF_BURST_SIZE 1
`define NVDLA_MCIF_BURST_SIZE_LOG2 0
`define NVDLA_NUM_DMA_READ_CLIENTS 7
`define NVDLA_NUM_DMA_WRITE_CLIENTS 3
`define PDP_SINGLE_LBUF_WIDTH 128
`define PDP_SINGLE_LBUF_DEPTH 14
`define NVDLA_VMOD_PRIMARY_BANDWIDTH 1
`define NVDLA_VMOD_SDP_MRDMA_OUTPUT_THROUGHPUT 1
`define NVDLA_VMOD_SDP_BRDMA_OUTPUT_THROUGHPUT 4
`define NVDLA_VMOD_SDP_NRDMA_OUTPUT_THROUGHPUT 0
`define NVDLA_VMOD_SDP_ERDMA_OUTPUT_THROUGHPUT 0
`define NVDLA_VMOD_CDP_RDMA_OUTPUT_THROUGHPUT_USE 1
`define NVDLA_VMOD_PDP_RDMA_OUTPUT_THROUGHPUT_USE 1
`define NVDLA_VMOD_SDP_MRDMA_OUTPUT_THROUGHPUT_USE 1
`define NVDLA_VMOD_SDP_BRDMA_OUTPUT_THROUGHPUT_USE 1
`define NVDLA_VMOD_SDP_NRDMA_OUTPUT_THROUGHPUT_USE 0
`define NVDLA_VMOD_SDP_ERDMA_OUTPUT_THROUGHPUT_USE 0
`define NVDLA_VMOD_CDP_RDMA_LATENCY_FIFO_DEPTH 8
`define NVDLA_VMOD_PDP_RDMA_LATENCY_FIFO_DEPTH 8
`define NVDLA_VMOD_SDP_MRDMA_LATENCY_FIFO_DEPTH 8
`define NVDLA_VMOD_SDP_BRDMA_LATENCY_FIFO_DEPTH 8
`define NVDLA_VMOD_SDP_NRDMA_LATENCY_FIFO_DEPTH 4
`define NVDLA_VMOD_SDP_ERDMA_LATENCY_FIFO_DEPTH 4
`define NVDLA_VMOD_DMA_LAT_FIFO_DEPTH_MAX 512
`define NVDLA_MAC_ATOMIC_C_SIZE_LOG2 3
`define NVDLA_MAC_ATOMIC_K_SIZE_LOG2 3
`define NVDLA_MAC_ATOMIC_K_SIZE_DIV2 4
`define NVDLA_CBUF_BANK_NUMBER_LOG2 5
`define NVDLA_CBUF_BANK_WIDTH_LOG2 3
`define NVDLA_CBUF_BANK_DEPTH_LOG2 9
`define NVDLA_CBUF_DEPTH_LOG2 14
`define NVDLA_CBUF_ENTRY_WIDTH 64
`define NVDLA_CBUF_WIDTH_LOG2 6
`define NVDLA_CBUF_WIDTH_MUL2_LOG2 7
`define NVDLA_BPE_LOG2 3
`define NVDLA_MAC_RESULT_WIDTH 19
`define NVDLA_CC_ATOMC_DIV_ATOMK 1
`define NVDLA_CACC_SDP_WIDTH 34
`define NVDLA_CACC_SDP_SINGLE_THROUGHPUT 32
`define NVDLA_CDMA_GRAIN_MAX_BIT 13