// Register NVDLA_CACC_S_STATUS_0
#define NVDLA_CACC_S_STATUS_0					32'h7000
#define NVDLA_CACC_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CACC_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CACC_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CACC_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CACC_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CACC_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CACC_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CACC_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CACC_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CACC_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CACC_S_POINTER_0
#define NVDLA_CACC_S_POINTER_0					32'h7004
#define NVDLA_CACC_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CACC_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CACC_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CACC_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CACC_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CACC_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CACC_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CACC_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CACC_D_OP_ENABLE_0
#define NVDLA_CACC_D_OP_ENABLE_0					32'h7008
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CACC_D_MISC_CFG_0
#define NVDLA_CACC_D_MISC_CFG_0					32'h700c
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2


// Register NVDLA_CACC_D_DATAOUT_SIZE_0_0
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0					32'h7010
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_RANGE			12:0
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_SIZE				13
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_RANGE			28:16
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_SIZE				13


// Register NVDLA_CACC_D_DATAOUT_SIZE_1_0
#define NVDLA_CACC_D_DATAOUT_SIZE_1_0					32'h7014
#define NVDLA_CACC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_RANGE			12:0
#define NVDLA_CACC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_SIZE				13


// Register NVDLA_CACC_D_DATAOUT_ADDR_0
#define NVDLA_CACC_D_DATAOUT_ADDR_0					32'h7018
#define NVDLA_CACC_D_DATAOUT_ADDR_0_DATAOUT_ADDR_RANGE			31:0
#define NVDLA_CACC_D_DATAOUT_ADDR_0_DATAOUT_ADDR_SIZE				32


// Register NVDLA_CACC_D_BATCH_NUMBER_0
#define NVDLA_CACC_D_BATCH_NUMBER_0					32'h701c
#define NVDLA_CACC_D_BATCH_NUMBER_0_BATCHES_RANGE			4:0
#define NVDLA_CACC_D_BATCH_NUMBER_0_BATCHES_SIZE				5


// Register NVDLA_CACC_D_LINE_STRIDE_0
#define NVDLA_CACC_D_LINE_STRIDE_0					32'h7020
#define NVDLA_CACC_D_LINE_STRIDE_0_LINE_STRIDE_RANGE			23:0
#define NVDLA_CACC_D_LINE_STRIDE_0_LINE_STRIDE_SIZE				24


// Register NVDLA_CACC_D_SURF_STRIDE_0
#define NVDLA_CACC_D_SURF_STRIDE_0					32'h7024
#define NVDLA_CACC_D_SURF_STRIDE_0_SURF_STRIDE_RANGE			23:0
#define NVDLA_CACC_D_SURF_STRIDE_0_SURF_STRIDE_SIZE				24


// Register NVDLA_CACC_D_DATAOUT_MAP_0
#define NVDLA_CACC_D_DATAOUT_MAP_0					32'h7028
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_RANGE			0:0
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_SIZE				1
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_FALSE			1'h0
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_TRUE			1'h1
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_RANGE			16:16
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_SIZE				1
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_FALSE			1'h0
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_TRUE			1'h1


// Register NVDLA_CACC_D_CLIP_CFG_0
#define NVDLA_CACC_D_CLIP_CFG_0					32'h702c
#define NVDLA_CACC_D_CLIP_CFG_0_CLIP_TRUNCATE_RANGE			4:0
#define NVDLA_CACC_D_CLIP_CFG_0_CLIP_TRUNCATE_SIZE				5


// Register NVDLA_CACC_D_OUT_SATURATION_0
#define NVDLA_CACC_D_OUT_SATURATION_0					32'h7030
#define NVDLA_CACC_D_OUT_SATURATION_0_SAT_COUNT_RANGE			31:0
#define NVDLA_CACC_D_OUT_SATURATION_0_SAT_COUNT_SIZE				32


// Register NVDLA_CACC_D_CYA_0
#define NVDLA_CACC_D_CYA_0					32'h7034
#define NVDLA_CACC_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CACC_D_CYA_0_CYA_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_CACC	32'h7000
