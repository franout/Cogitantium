// Register NVDLA_PDP_S_STATUS_0
#define NVDLA_PDP_S_STATUS_0					32'hb000
#define NVDLA_PDP_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_PDP_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_PDP_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_PDP_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_PDP_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_PDP_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_PDP_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_PDP_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_PDP_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_PDP_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_PDP_S_POINTER_0
#define NVDLA_PDP_S_POINTER_0					32'hb004
#define NVDLA_PDP_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_PDP_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_PDP_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_PDP_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_PDP_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_PDP_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_PDP_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_PDP_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_PDP_D_OP_ENABLE_0
#define NVDLA_PDP_D_OP_ENABLE_0					32'hb008
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0
#define NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0					32'hb00c
#define NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0
#define NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0					32'hb010
#define NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0
#define NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0					32'hb014
#define NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0
#define NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0					32'hb018
#define NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0_CUBE_OUT_WIDTH_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0_CUBE_OUT_WIDTH_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0
#define NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0					32'hb01c
#define NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0_CUBE_OUT_HEIGHT_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0_CUBE_OUT_HEIGHT_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0
#define NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0					32'hb020
#define NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0_CUBE_OUT_CHANNEL_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0_CUBE_OUT_CHANNEL_SIZE				13


// Register NVDLA_PDP_D_OPERATION_MODE_CFG_0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0					32'hb024
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_RANGE			1:0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_SIZE				2
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_POOLING_METHOD_AVERAGE			2'h0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_POOLING_METHOD_MAX			2'h1
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_POOLING_METHOD_MIN			2'h2
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_RANGE			4:4
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_SIZE				1
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_ON_FLYING			1'h0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_OFF_FLYING			1'h1
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_SPLIT_NUM_RANGE			15:8
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_SPLIT_NUM_SIZE				8


// Register NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0					32'hb028
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_RANGE			0:0
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_SIZE				1
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_DISABLE			1'h0
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_ENABLE			1'h1


// Register NVDLA_PDP_D_PARTIAL_WIDTH_IN_0
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0					32'hb02c
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_RANGE			9:0
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_RANGE			19:10
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_RANGE			29:20
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_SIZE				10


// Register NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0					32'hb030
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_FIRST_RANGE			9:0
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_FIRST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_LAST_RANGE			19:10
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_LAST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_MID_RANGE			29:20
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_MID_SIZE				10


// Register NVDLA_PDP_D_POOLING_KERNEL_CFG_0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0					32'hb034
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_RANGE			3:0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_SIZE				4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_1			4'h0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_2			4'h1
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_3			4'h2
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_4			4'h3
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_5			4'h4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_6			4'h5
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_7			4'h6
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_8			4'h7
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_RANGE			11:8
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_SIZE				4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_1			4'h0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_2			4'h1
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_3			4'h2
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_4			4'h3
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_5			4'h4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_6			4'h5
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_7			4'h6
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_8			4'h7
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_RANGE			19:16
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_SIZE				4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_HEIGHT_RANGE			23:20
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_HEIGHT_SIZE				4


// Register NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0
#define NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0					32'hb038
#define NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0_RECIP_KERNEL_WIDTH_RANGE			16:0
#define NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0_RECIP_KERNEL_WIDTH_SIZE				17


// Register NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0
#define NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0					32'hb03c
#define NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0_RECIP_KERNEL_HEIGHT_RANGE			16:0
#define NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0_RECIP_KERNEL_HEIGHT_SIZE				17


// Register NVDLA_PDP_D_POOLING_PADDING_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0					32'hb040
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_LEFT_RANGE			2:0
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_LEFT_SIZE				3
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_TOP_RANGE			6:4
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_TOP_SIZE				3
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_RIGHT_RANGE			10:8
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_RIGHT_SIZE				3
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_BOTTOM_RANGE			14:12
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_BOTTOM_SIZE				3


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0					32'hb044
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0_PAD_VALUE_1X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0_PAD_VALUE_1X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0					32'hb048
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0_PAD_VALUE_2X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0_PAD_VALUE_2X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0					32'hb04c
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0_PAD_VALUE_3X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0_PAD_VALUE_3X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0					32'hb050
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0_PAD_VALUE_4X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0_PAD_VALUE_4X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0					32'hb054
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0_PAD_VALUE_5X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0_PAD_VALUE_5X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0					32'hb058
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0_PAD_VALUE_6X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0_PAD_VALUE_6X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0					32'hb05c
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0_PAD_VALUE_7X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0_PAD_VALUE_7X_SIZE				19


// Register NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0					32'hb060
#define NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0					32'hb064
#define NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_PDP_D_SRC_LINE_STRIDE_0
#define NVDLA_PDP_D_SRC_LINE_STRIDE_0					32'hb068
#define NVDLA_PDP_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_SRC_SURFACE_STRIDE_0
#define NVDLA_PDP_D_SRC_SURFACE_STRIDE_0					32'hb06c
#define NVDLA_PDP_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_DST_BASE_ADDR_LOW_0
#define NVDLA_PDP_D_DST_BASE_ADDR_LOW_0					32'hb070
#define NVDLA_PDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_PDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0
#define NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0					32'hb074
#define NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_PDP_D_DST_LINE_STRIDE_0
#define NVDLA_PDP_D_DST_LINE_STRIDE_0					32'hb078
#define NVDLA_PDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_DST_SURFACE_STRIDE_0
#define NVDLA_PDP_D_DST_SURFACE_STRIDE_0					32'hb07c
#define NVDLA_PDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_DST_RAM_CFG_0
#define NVDLA_PDP_D_DST_RAM_CFG_0					32'hb080
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_RANGE			0:0
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_SIZE				1
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_CV			1'h0
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_MC			1'h1


// Register NVDLA_PDP_D_DATA_FORMAT_0
#define NVDLA_PDP_D_DATA_FORMAT_0					32'hb084
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_RANGE			1:0
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_SIZE				2
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_INT8			2'h0
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_INT16			2'h1
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_FP16			2'h2


// Register NVDLA_PDP_D_INF_INPUT_NUM_0
#define NVDLA_PDP_D_INF_INPUT_NUM_0					32'hb088
#define NVDLA_PDP_D_INF_INPUT_NUM_0_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_PDP_D_INF_INPUT_NUM_0_INF_INPUT_NUM_SIZE				32


// Register NVDLA_PDP_D_NAN_INPUT_NUM_0
#define NVDLA_PDP_D_NAN_INPUT_NUM_0					32'hb08c
#define NVDLA_PDP_D_NAN_INPUT_NUM_0_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_PDP_D_NAN_INPUT_NUM_0_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_PDP_D_NAN_OUTPUT_NUM_0
#define NVDLA_PDP_D_NAN_OUTPUT_NUM_0					32'hb090
#define NVDLA_PDP_D_NAN_OUTPUT_NUM_0_NAN_OUTPUT_NUM_RANGE			31:0
#define NVDLA_PDP_D_NAN_OUTPUT_NUM_0_NAN_OUTPUT_NUM_SIZE				32


// Register NVDLA_PDP_D_PERF_ENABLE_0
#define NVDLA_PDP_D_PERF_ENABLE_0					32'hb094
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_SIZE				1
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_DISABLE			1'h0
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_ENABLE			1'h1


// Register NVDLA_PDP_D_PERF_WRITE_STALL_0
#define NVDLA_PDP_D_PERF_WRITE_STALL_0					32'hb098
#define NVDLA_PDP_D_PERF_WRITE_STALL_0_PERF_WRITE_STALL_RANGE			31:0
#define NVDLA_PDP_D_PERF_WRITE_STALL_0_PERF_WRITE_STALL_SIZE				32


// Register NVDLA_PDP_D_CYA_0
#define NVDLA_PDP_D_CYA_0					32'hb09c
#define NVDLA_PDP_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_PDP_D_CYA_0_CYA_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_PDP	32'hb000
