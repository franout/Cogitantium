

module filter_and_select (
input a
);


assign a=0;






endmodule