`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TzqTWzVLLXocOg3up6rNft4bohjJcXyx5Czce07G9z8MNQ+t4/kAN+nY1jVADeFtec4dkdZh45H7
dpcDQQdQTw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z3AIpLDjUuaEQmH82FVi2zLywElh7iOAf1iLbsH/YfB5BOyx+3wfmVCJ6Zjar0dfRtQcv0eQfDcu
bSYBTssSuSkuCYCY0rBpM+Xkdyc7/Xpr3LQA/00f0DEGwnxc4k0YsovbPLFcIRhvP6FJgb/UGXjN
GeLE3Nuj/DFsjPWAUWA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
seLkBZQbnIZh8mBM0T8s4G+scEHnQv3scD/jzq5LdHSnBvJ7KWwKEYrQa5ly3MWqO8Vb8VGHVung
MRPCKAbHQm2xgx/Uvhde0GLcfxIVTgX3kJm/0+Bv2q76aFQujYtAgg7uFAAwhyAkkfnHJ/A/aBIW
xh9lJdgtdUmQAT6Z6KA8XqCpsm/DWgKArIz634L2J0CrcyCo46iU6hGrAn45XPYZZBox9ahEUs6r
5mKy0gW0d0uleyI0ZrTMugAxjdGKCjei/AExoShQrKErb8/wnmsGgiTVh28z4pEFqLq+SZuHd2sv
jeLtUGm9TJ9bxz5LprsO5WCPvzdNC3OYYbnpgw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DiPRLFQlcSB/5cG25z0ajZZB3DoqPLpKoD0KRMKxlyW4WsaFtkBrkokE9RoW2RgsVy/ZaoiS/E7R
jJu4KreD9pe8InxBB7i9EvvgY0v4ddCszu6rnbqeYPCZz6IbdT+ymjZWCr36E0XT66t5NuRpERbP
df/Q7vjXkz48MiNmr0HCKN93gTwJDzxzOFLPlKJlxV/KmdZ91J7J9T7g5u/aIqPzQE6e2+gEAtN/
Iur9tKgBhdlZ8rNYJwBZTKs/cn2fp3TNG6eYzzw/goWVr55yC48vjFpXrKH0QX5HIlk1VIS+P5Jo
Ovttt6MLNHbEBD8FH0DnWdF9nKLTNQtZ/AE6Ng==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VQJvMecUTSyfwFPpZYbnyS8ZLP9HSCVo0KZIrrWWgmtNSfxCEVxc1wJA9rQctCqMtTSrapXwP1TL
imlvt4vq+5WfFdAzpSS+XRfcRciD1B/o96Brzbf2d6h2S8/Q2ZQbUolX8p/4kLawMrL84Mtncm9C
4bIrtZmPOMxCa4HtYP/go4c7SJpV2gTOGY7zY4SXPIA2VXGMDF47OruyLpiXgEWfJXR64iZO2f9g
R+v1qeda455LtzSv7VaEnbTNJLcTsZksj/jzZrjJKXFFZ5oBftTJpoA037hbCJPEti6nXeqO8kf4
dJPK/ghG+jCFoeUk8LYz/L8xKEoOzOrCjmYsCg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C/BT22ARqkup8t9IdChI5dvaOZ9kZM4efppnEoskwNGXu/0HBwEKIB4bPBAXgoBFlTJQgAC4eXI0
MnSH47MSH4Btm4q7hJFjTef3V1YbSOJma1DYl9f4GGud6Mw3AiPAacUsu2LRpCvvaIXx3o4nIOFH
p90yAimODI6d7n3gdSo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZV/QKk3FV4ZMZVfsG/Zb/2t/+6f8be2xqgHelh3OLiRzE963in81thjQvazEc5zc1n4owsRx2ORb
K9UNCgfm8uzAjqZI0Know2dOFLKV4yifU15QXwPabJad8KkfNxch8e42iWkDU1gM3pX9TZU2M/B7
W5EjY212YGfIOUSbz4t3AEv+s6mIe8+Pj3rEp0TJi0i3qPsoTlcfOYWGrMdedLLbgGCk9g+X9sCF
ipC6cYcKQUt6O5BHVpjngy2zzVQvWDTAIWRjQURcKGK7/mfaw+87vhuQxxeTq0Uduc6NZOFXy7hf
zCHbqhG86f7kX+A+VUQCO7ZEXtiIDlYbJy+ZWg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JnlR9DnVIpJP1LXCzYrM6mdoqOotbn9RJxUMSn1U1dN+qeyzM1JLPN3WvXAzafxhzQfg/b2OXS0b
VljW/hZBWuyGad8AOSTqi68oMMaZmPtGJn8WbGsVdpCeHHDkeXU4+qtlc6w9LYzICJuZrYZrAGAw
bT0PjT0r0lgHw0FNdlXxlfOCYwl31LKHexS9ZtJjMYI4wO09BS9OLEjzaWQT92IcBA6IhcAKk4lv
+KJ9Hditqjb0QuKzSPTcREM0V4QSTXJP0lW81M7G/XEVwTx82QoTrk8AhHQhJFLPRmIrfoF7DTc9
sOhtub+eZJMrCoTjpWVjYj01gaq5H4jUlDblXw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
djIblLtuL8PEzD4uw9iktIXCVe6CopDcg8vmC/R51+cARhYEblBMInp815RGUjc6Tw+zQYDB14uC
ao8/VmgAEyxuL09SwHN5S0FzpvKu5UtLaPdVABYYoLBj49G3fFB7WAvZ4aGo84hQSI5mXBVhWZg+
fl6d9Vkbo/mbi1+K8s458g7FLRp+kIGXyn6iYGPTzNaClivFGHCt66wSvtOyPqK034GkpgShHs1+
fUZyDLQZvifa68lPnA0yIipgEnG9UWMsNW4GDgOJaC4JgGjj1VUKh6Lh6Iyr/hje8nbh5O0oyhGm
59SDbh40qDfaRMKwcfzgFhdK9w23qsIiyNofUy8o8C41r1XU6HJ02dd+Gxi/wT5QhNprk7QTBebO
rv4rjG0YFS8QEGCi5p+zbN9oLcF3pNUWaHog2lFJcZiyJA2VuHWxcQ0XfY6JZBeVOyj5LS6o67zF
F3SjEet8q7lv9Ha3k87YF5L1F7D1dG6AAfU9qKVYW+k92x2f42aYunDipwH5EKA3Ci3r8KA8UJb4
bDj7dr/e9zAyBRoiwXFGzAqkYM1dKN1y68wjxA4jE3otCnxqpjZRGXftyurZ5Ku/40Q34tsWL3Tk
03klQLm5+szP7bvGWQOv2xG3ltEx6ygOV8/TQzBjJF/QykgSahmxlg9SnRpxDebmdCKwKSzn/jRh
1+y8nKsOddQElZ2A+1oX+CXubv7uLdcEC1oi9dhOGYwutEFdH8tZ5slIOZaowxwlvdkFAVQlRnx1
HnirNv6H5mThCKmlArFl6fuALstSCWcuMNm+O7bYZJ4sL2TVN4qD7S6LPc7+2JdwgSFc8FEb5NrQ
vIBkn7FK2HLFlLMHoHeqY0B9W4t0dfkaZniCqY1ULgqst3iUIKM8GKgcdM1hnL8R5DrLVUKYa1XA
lGbEJr8JtUXa2k3Ccye5ijbWHBUHvqG3LIVPwHR/ltGvTwwNWleZdhFmWJ7LuKvrBxv1e+7Rh5F5
o7UEj/dPPalRGLjadwzwPoxFg5xbmKabAq01O7M9VzWsY03fPxQ31nYWxJc0P4A5YdwdAosbJAhP
LdH51jWLkaXVMrTzM3nJjq25y1zSUrvivyqA8v1K+1Ph3/W5GIVxhy4QUoyJ3nyDT2n/AJVyY/vg
uYTR2M+7JNyap0YHprvffPJoN1w94kh3/VuesOg2/jA8gwA7CinTdU9ScvJ4e7vxNC1jLxodM8S9
S8u7O3yzM8/BbV/Bhb5vzRv2+NSK7iaWZWrn6bgvoqGRywlyEP6rDU+/9FuqKk6nOWHRGfa0JT+q
4yckeaNEE9yAsToUC/NaW5gATYqcbL2337cbpxnvyMSJOvKtGX2dOlZ7PDaNxSofKOzeJXkU62g4
WFO5qUTYb5Fj/Ctv7GBr7HzWhDhsoJ+ai7f/wFzMqi3SAcg81ZH8/4ZkwyNde42S1q98ioHYCltj
MJHbtZUzg2g8LOz/GH4h6E7Jm73xES+ejxs0zltdPkA0CjKHXPJ/d3q1FUZ78aw3EnnGiWuVaQCk
97iykThvLkeFytbBADuPMGIXP5siTtIhYFzuGQ7SrxWfltSHW+lPjgDFOmCSpeSMDeIHgy38L2ap
SuOMQ8PBs5dVXXYV7p9+89U4WwhLkAz07/K/dDb66ulm5e0rksuYU+xXGs3sDQzXQdmcXfxBcGg4
9fK9VBLNbmH6zF5Psu1YboT7kOMDRgHvxyHgn6TmfZtBLgKpdt/8vf31ue7Hg5gGrosm2RGEwpro
RzDXt58AbPUNlwVxtdeOMd6loJiGxK/GD8lDmDaY3/uOTr+wPsh0szouC+utprcvNawsfOVYRPW1
hJD7UxDvvfvruPEfGHpYxK99G1g++/atLWwQnvLYZTMf3KKx4SUb4MmjNjuiXCm0PpsCvxOsagti
1YQbzX5WL7u875NMWeFMD5ViHDORSDvRMqKy1tSw9bp2CW/d2tcRXENyo8P/4c7RG6/ccxs3wv0u
CCbuvYoJARnwEeJkSvIAMUvN17KFNyBnPylo8Lr/xvvIUL1mljzTTU1A79zUi4A4IvsMyqgLm2vJ
n7eGgDYXVs8hhUMZJIMk++DhCIeLLOQpvQNHHLRwKn8rv/AU3NFa1XEmYj8Ph2wFZRTyDeGomEKn
Wt/VlD+MlDc39aFYxHxto8Ee5/7pCnZwc2iOiigdcIrMuF2+9dUs91A7gCome6a6YKGnrYgRzJsl
/s53L3AAT783s+LSKFZXtsxIR4zG+irvXWd4ZJz8823AdQoRAwN+8uWa/Nu2yHcKn9xGxctzNWaP
cLIIw96Ap+kDseoZuD1inhGVTivRFqY6FjakWuoemzVupf5iJ67IQUrUnLhUop/351s28sk10Ud0
jJ2zmoHzk6RN6+BnNUTWrOFDA8oJLIPyKWgpWy/PFJxyhj/flaaX9w2MJaVYrxX8dAz0m5tYNaba
n3kicOjXTsgXm/AIG/1eHSB/9h8rCK5262ah1TVCmYrP+ad0+CgPbgTYleL6URKLH+vN9TPGUtoK
ZdnkuJLv/XU+zGberELu5mwuEqlD+kxPLDfUb7VCfSq1PGFwPzePoZrcS1gOzMgS+6ekWWJodgRA
CU9eKsrmyU4BFZ8MNs3mSwcfuRdV0dmAHxZLvFeVY8n9CT4oWbOhMwqY1WzX/tQM7sWwtZ6TsWz9
nlxRn3Sg/KRqeg2Cc5oxvOuTE3LFdrAgHDnggXGJ/j61oCOIi1nY3lthQMrJwCOJsX5CTjDUAPaU
D5NcchytUPtjR2Npn90e2Y9K86DUJyYGUlt2nFPmIU8arPbcjLfHUyjir0xNh6HkN2z7VPg6etbk
qWXCuxgFbDjHeHeu/Jc9q0jwcu4KSD8zZTkdxhENs11Xi3FAiCJFsfLQE/cuQ6Zx//jVEjgZ6qRf
6qOGmtlTyeB8jTdygF8LSSp2LZArImSX0jX7SFUxNkQ8FMpDFUauzHToslPj7n9xCcV+TQHMkaTt
aebync3QD3ZPfhvv9Sww9AxMmaFwf7sctSMmPnGX8njyKkzvT99CXHkF//W9121Q/XeZNzTvSUmA
kckDQ5gAovU4ydAIr/v/S97We0rjv/Ki5jG/rXQTnYyq5Qllv0gVQuMDm2R4JQEgd2hh3T47vOdt
NqoRFCLMEUoZUtlG8SQPRv59KAV2SEmhPctny+i7xuYoekz5XyJsfkfC+ckHvB6R48aoosh0H7Nf
qzTaM5RdEvdzjO8x5AZiljEcnjQl8oD7zc0tEp+7UMdtYonLJOIsegRsGgG9JM0DsMLAj528Gtek
CYLiFIjMNi4VhLZnxavAuESmwi0Gs0HKmpIEV25aJZoL6lvjN0meT+Nm3AyHBYMH67eo91CeGtbF
UZSieZ6+CWCOvfz2wi4jIF4luUyNO+dyoYSyHV19tXuaWaWmR3u59k2OgIxvJhx86ZUDJYgD9Tty
HFSm7zipERLk4cLYe7FXhrb2KaxEJlxG71iz+YlR3ViZIILZWK1yp24MrbnOUdBMdB2Uy9vEampq
vUg87UDtsuzobravNrjAJEScfinpUEV2cdQWtFkLcRsmOUFUef+Uz8catgvVAyg5Q9aeU/qiqneo
/FW/UlGZH4xiYnPgd0kN4tEXcKx0Cvp/SE7X+2/ttF9LXaSgISN5OmmLzrD3eUMHaOEbzJUUtvim
FQNR2db49yjkN7Hp5Tk5tP3M1Gw8VyaUspUSx1oQGLy/ACr81C0HqkbI4J1QyyNAAmWWboqYiMRU
etOEeTFlxJo44h7nH78pQn1kGGZQAE4Sgl5qncSIAWOmPR+AarG+taDPNIaK/5t9+M23hdKj0M4G
VSiX2dmKyqkmChll0YgIptSRP91FqMmu8iyaelmMoycTwQdQfK2XClZlJTDqmybLVe/9hqLAJDGA
d4hDTMdOwW9SwzeO9r/DjsAeUhLOlXJVyLHPLHuC3aeb3rf9Y259wPb8d4Ao4U5zwzu3fNvjd3jU
Qwp0eZaoBJNA0N262+68sDfRKll1mOubDzBz2MOAf2AIpsUhomtQ9RuHt9f/PobLH70v+oGYJdH5
H5FthrE+bSEEIFvMfq4Hxb2/PrVuPKByhmis3QBNpr2CbzpdsiqF4glicsCFh620FhQUONWPAPG0
z/CoRa9FFj/b3Vb+dz0w4j+LokZvxCjuP0Eyge/Rkw8jo05wHVonG5C/KUK+sStRXi1cAsjtvFUf
t+gkvGoygPNRmLcTYNGcW5FTR7RBIJY5cYX2JQVYJNYJNrLr4hf+rvAqwimB659kNsc7Fu0BJgC4
0kTxfPgZwoq1KOq+DTMGTDSSJBAhGCGfIVgfwfq3bNXzsBhbK2Iv7BLosExRZ7/oMO3GRghAOZtV
670G4GMPqoQMmQnsm6OxQQzuRxX3QfF+qvLm/Cs01YsUlLbe4xTzFQg8FfMWyD7atk/YrQ7ZpSVo
SD9kjgOyUAdxz2PVDh8c0ssLugx1JLc9uXt4RH6Cdyh1dRVKBanJ3fBSGh0rL5Ph1bI3ukdlVrBG
FdWKzA99huv4dERQN2ilZVeLB+xnoUxPv6ht95S+MCUczDP2hjcnt9BZz3LlbPNYx4GrSnrzQZB/
+SLsjdCb+zaa2o7HsUJmwTTdwA5NRB6451yJkpcj2LRG1DWfUdGxtWIgbK91da3fNKuzgXN6p/C0
vTWiCvOt1T4g93ZTvVj62y1hnE+8OtLhw6yGcuNBMLi7rJxEKZBrK37TNgmqdtsPZiCBEsB+6Uie
CCxNCIivatplxYdRlvEu4Wzn79cQ4Ii1ZqAZOnKuGZUOSlw+jGh5nqZPI0CzY7BlYVH9+95tH+rM
N8znI5Ev3CwTyf/z0/gUyWnUbaIC8u2N+kMi+9iR+YPjCUVkCMYvBG/pnMVVbVzYEx2GkvQ65w3n
2jVFeke2Vy7P5n2D4aNEejGiadVbJ4wk7LTUxGr48bNpP8/fQh4CJYPiMLCkvl1EJk21VBazF0IX
SWYPpUIDEXMLqLiP4eJPIIgHiE65+aXTqnO2T6/nVyF7l21USU/pOLY7zXhqozcOC1dwXfcJP6xd
cCPiBV/gin6/NpwZlAlfcE5T2ktPqJlYuOgF+iRmAbPbPMR8kF9FVOF9xPbhZYNQAPnXHbcRyW2b
wb0qoq09ScMbmZRdfx6WHS/GrTBpWKAePspZUT2hdoh/Qe1h4phFxMg5cOCWt9ZuJSmAosSaB4l3
lRLaoLuIaowFRlg1lXTcRUg1K/Ni/tC6Dp4cBT2BwfAv/qpDpkyyt/UiDzIRI+wkZcJBufjMhIB7
l4wuRA64nkqBnUAKh/l3eR0pVVsJ8JVYBD4rZfBQ0a1SexCK+HvKvkXOyDR5Fu8m/RfsdKESnjRa
UQAHzIZ09QKt5jB3ljuj3RyF0wk0vlJFipG3TAe6X4cfLOQvt3Pd9eWh7e4fm/MQ7UerxSthGnWz
OrFeQcnhJsYzm0CROSH8niKmoxCjnGUTiA6azbUAU4E+GnEI/7Ijtt8BRdZc1wM1Dp3wvOEzGpOv
hjDgakMVDggirnK5bbaRL+3LCAeNRSN7xEPFEhdUBj/C6hSaaUlLiKJeCRerVw2y2fSGbfGkym3Y
qKVhJ7wk6Y5HSW1+dZY64hEGK0ZxWQV9eg5aGzTlOJRzucGrj8DEnZwfEVKVF79QYha26d3UMFtR
kaDr624bt1kiH+OEiKV9Qaly511T1iIr0G06pIDhJiaSfW1UkWivvrh2Gwhv9HRblcrbnPvLjuNk
phqCaF4hWXrGKSRV7YW6oWc193atQBXw3elFhGwvRK0vMMzMTzFNKjm71wTPzXqEAbjq5quO5VLG
gMkzmSt2NuEoEryhioyKLgFvqDNmuSRnURVs9z9YjiRroeuEpl0FWAUA0nvio8GJPWTWbYxexZO+
EyfxtfH8RHpeYRPdPPTKhnbNg5QtGNhz1KfD8jQ8S/Or8y/EwMm0ctRnjmPaQgoi/cCVJbeif4nF
JpHOjpk8Vz6uov2bku5kY3xER8Qgxy6BSE1BaSIR3CA7bQFNwEiq0oD5VQYnJD/xyIfjiZj7OpEG
+kAsrBePF3CZGPsAWwZj2np50ICFtkrkLb/CxN/cDPdPSSCumE0M6Pb0rexQMqH59NG+Vv7jeaE2
Ew2FBjXAmiwPPGpJsjdpuG++DAzZQTLEasTP8KAYTIfO/uyhgda/pq434LMNKrIw6/GSTE2t3t6e
LazEhO/0ThebGATPf2EfYqfa3zsXPhGUEfugoiNSrUXr3vyeF5RLlSo1WWpeem1JRcfOu9uOltLK
1xhArZHt+rA/L2/d23St8bav8OhwvmPD8jn8pfVhkfpRUgOK3iRFm+j6a3ME4YNJd0oCl6JakRvE
fayKEBOsjWbn4AgdGd0Hu8xDVFIE7tgeMTVwHoES1GWSL7ZOUe3Rwdl57hiUqo5sk1wQEkMxZdpC
/VKVBH0IH18oqQ1b4eIy7qobTF4WS7p0CmAq5yvZhu50t/MNKnMWXfMYRohePLF8C54jAb2RoPhV
8uOni9r7lRR/5xy33GlbuGbsO2WBPlJGukwRm/NkMpsiFBH/qXnuZQq60Hqe7PgBWhyl9seAhtnb
JbrP4WvBVuOtmiNl1AxyH/6T/gHmyy4kTb6cyzhyGm2HIl2p9pJwEpIMqoJFJhAaIIoofdLdqYUw
tkJKurnmQ/D/l7LCGU0oDp9iEMX6CM7jXUPpMVb3hjISgk6fH57JcRhxs7C/hdniovanvED73bLa
XP8g9RfLqn2Dsn5fBGB/oDIJhL+DjLqK+r5zruqBrkD3G40qw2rzn1+jkFlzz/zbCWhpQW3ouSXV
P6joSRe4tpP9qzT4/sw5IjGlHOWZ+hna5hVMScWlkqFoEJRLrJtclTsZg2wHtwsq+WBvbnfmAezQ
go1Wc1Zb/WcaA84RFW8ZK+rwFEag885zDifaSlHdeWUDObHYAhnv4IG67k96BtT/lz/4/COeaYeB
apL881sA60dUfKpE0qKBmJRpgH6XSPeGI0eAOJL12OLRGrA0bGxehGriDSxRrEV6h/W+IpHRZOlM
8BZsMtNG+bgGxotOSwksr5LDcV4nK80QdCTFVLU8lJjDVdR6vjAwdGOmuZsxB5ehTfb+QaOLycVb
5Z1q7Ec+1Ka/xVSyGRf6lyi+htPl2hh8WQMd0OO888sHiBeSM1HPkHQVNvEi18vfwyYpQtZqHduR
Li+aIvIGZFcLPD9utHeuxLO7GH66tgdx4pI0qFmVwllWnWOvcxQNgRIjIRCHp/DOI2fT8sIzwISd
szEQuU0MO0SmFEZlTdiooJ7NTJZxN/qns8/iiz8c7y74Wh9TF8+fzkOcFNSUMzaQmksKmNjrpm/A
dysFbRaW2DUrVyWY4WBdVKhpWE+kn0+8D/O6XI6YRkivVWM/hlWqAKzK69XS6ZkZFd0PUrjKiaBV
oPJ+SzF8Xp1TNd6U7NLCOY7CI4oDCeH1tznVSOgwey8JKBHkuuhk+HPgRxyx2I2XbA5obFuVkVMe
UT7NOAiAWBJ0okLrx47bNhyqIJq+EBl1CB6VECxL9SnUqnHEDd9XBkiCBANzboLoNLPjw7erZSUa
Ru4tqustuMEWZVL8VuRazyrgWyzapOR9CFqgiXw0cRBuB2VpeqjRFyfn3tjY1JMbukrgO148N7wB
xOcWOt6P0QSafCLQpgw+P01hLpPuYGvQQyrm92mpUJNnZxqo8oevMx3VAB3RpgRZ5+sxHxuocecW
XTwzju4lFSiEyOdG7B//6tWVLJxA93RL340wnJj6SbPzmSn3UnLlbbfERfeLpnzW3HKycgQ6QORk
TKb134V3u7GQPcPkgduOipp/ePvHPLQHJIAT0HjTjYvzlKlBNBFvBIFyl3TimFic2/fI9FD6tw4Q
jKyqhYm/Sq3PoNYyAjdc/kT5VaFA9h+rwARnskPnp7+HAgCRD+7szo2WuOEuflmYetEEdeUTERXe
fMNk3sWr+L5RLLgD7Za9PWzLEOGGt0fVaRA12LSVhLcVjIFxwHbI5kjkocu5OJX8QulgZSgNLQMG
K15Ra8NFpElnT6vfe/jaMYThicE55KJ0Tg9+ozbusAEGxVWH80KcDiRJyOTj57tnOZABdu1/q1mz
kx4aMMgteeUOnou3WP4ellWLXinc/scokPGtNVDrrY7xOoQKx5YFXM5d04yvGK3WQdHVzgFcmwFl
ml5VdxqIUs+/ZcPBtw1vW6MryklOf3TDuwgw65JFWxaggc9edZU/svzjpWomAilnkpttc1y8stq9
hCIWgf8bx1anQzWyMtGDnMIrJBekYvlydytvlYd3cFiy/CV07qtx3n9UqC9+SY3CO/PR0xUEB4aC
jgev6CNeKUgHny25eZZcw6ppfOSHEzxS8gIKvkCvTlXYULbEhkSw4qYAw03vqOY+I+KVw/x98RhD
zKDccKv+3CSqDQDSe/4uhh+uQrsZRXmgZcjJTrDyf8HOqrkD3r+qzOhx27iL239lv8MtLKBsIWBq
0njqkGA1iF3onHWSGIHY1uLKOqM8ONWV86SNJxCDVFOV1GxfWIiBDVCzMqCs855MaUbyWgHXZ0nc
8B4xrDh8p7tK7a2jqVwU5z7/V20wPh3JqM6yGevulYPqbWX80AHjQjngvK4dSnLv27UKBI+N1p5a
Fvj2Bn3Tedda7pKET1JO+jI/h/GdK3OYdOTKanUjzPsPEhMXiQF63MVwmAqg8q8dLy+lot3de4Bg
Kx7xx3YfnI0pOeaChOjaDyoKwHn2y8UDX/kR3a72xdQCD8uJg+X8CagjPOPlDEXD46pbwcb+ox6O
uyPTNbmKlW0Fi7edEIUvbDgY93UVCCN54ErRDpHr9R/6lr7wMtYCMVTdPw62SXC7Z3GPLbOuuRto
hREt5va5vCWMGNCMFLP6HTovWH4l/K8MFeBaWkNAqXuOaN0g1L6B3sAgKhkzyYj1m6jnr+Vp2Hyz
89x1FwcLo6A9oQ4/eLtN85Xb55fzL8/PfxrAr+iD5O9L1N/AmNuAnjhsxFXKaVJlLqFqj+LC6SWS
mUg9nZ/f5RiP0C0jENO9U4rsfCAaDYG/Nbanl72eMtEnCgYeAZim54fsy2ZJKebOvlkQuj8WlnXk
8LyyATnbLb7NYyH5efKnuURq2bqIAVxPqrPcFDN3kP7zf6PTInQnwpjqzuAnOCXnv1/tOAXTYI8q
e1GHsCU7spfQq/2xERBX6TGU9hJs+MluJwuNFAzDR6pN2s72F4ql4AwKa8476pDglF5l3jXCn0xn
RsWmPUoNdseM7bsJS1PkoXeomaKo6zzgWMQbABDw5dRQ8TqWDG543SfWsONHIPZCexPW9gHpWskb
6UxdTNwM2QA/hQCL8MdykaX8DfZMjD4DAXdk/MBKysGqTj8dxRX+eXCt6UiXnzTkk2irPad+H3F8
r+XyfGece0FP+cMuoCeF9046l3ORXS3P+lAwV4AZE5KY+nEwPgmcM9bHCKVAzT7KMXGF+QzppsR/
93C4JiaOi1Psku/xNN/sToxDp8aJXcC1JVMdKm1TkrYKsc5SVbqAa0fXNEqLFaFuu+SoBWqIP5Yq
V05pYsb8dN4/je3T35X79Gz88dPUSAIyKYAxmyz7GI6bJ5Av83kVjgVBIGUo/d0sZ8snNJufm5Zn
In6yULz4/2+h910cLtTQ8uvONNAK9ZjzpmHu3ctshzVNzz9Th774ZnAB32fCjHFZm5BkydL8VFGC
6ZcvOP+74zPRAqtd/sqZJ2HWLmVBPl0bjluWvA8CoYVe0gvDrOUXH0qvB9R5yLJ+SZqrof5fpkZ0
hLvf+1MK9sB0NHWbAuH/+iMm/wNmlQvXZqGi/BU0R+Dde3VnI3htGykhmxEeLFHzU6k9m5QrT3dw
Dbw2yv4KPNZfGSyPjvTFPGsRKHmRCEqhs3H+d/VDqxclAPomsNBpyHrqgqOZTGataH+AorUsLh93
b5Lt1DH2X8o7B/c4kSze0uWkwvUeVqQGSutzImWm/V5pirfgXFM/By0x9sXezI0MKgd9UhB0nmr3
ifCAvp1yhw/YyQlxF1ptK1+8G8qhgRe9rfaLcP4K76nfRucxeae0vi/i1KWt5Imk8+ix5jVfJF5X
qjzLW5D3/auT3nkHx82vmedf1dd9bxTgoBybfP7Nk12UuiDR4makZVB62rBKNV45+XQD4XB2Xgu8
30v/dl8eYVg7I2w2dNLMwC2vWVHWaOLHb1hbQnLYb9stwkUwIzeIlvZWRtK5T+/cGmGLJnITY9ps
hkIuRCeEay6yg6AO14dD/yOXmvfZgXp9TfZj6djKJ1ZyulpiyJ3fHMQgBw8FKpJ3KhsKN2DpE2/y
ehEw6JQdlCTOAkCPWbqr2HILXi1XCxfoctaVv+fkNaneXV8qJ5Rjp4ZcjaGB5imx8bLXPN8TWUfc
/TdH5+t8Oy70U5QuaRD6vevZgUXO8wbx1l863aEftLpFrHFSNe9BNug69SzIrWzjxQdyU6fytiWc
olMCpX6kl9UeqYyW1OW+KJmhB+/EJyu7/lYIeawOeTneOSVlc6YGoGRSnQZD6E4VXr9fpky6EhAt
q4F8zDNNVzgOHYfD1m/ycbcz819LV4O7E3b80ZWGT2UB89dIHTyHM52CbraN4cNQFCfvPVGbOXiZ
AJpF54ZTjDjLAS/aE9ZpafqukkH2HAfuan+KzQPlZvSjRkCa9Zp8w/v+yJM2IeXorxogrNHBSVl2
EysjGy5uIZ8nlmgCRGpIq/cSCysYi9w/Tcht/nnBnv+nopLUBdwWVhAruEg1p8cLf0969Bf3cNeL
SFThOnOzYyqeeuatH/7SjtETIVcwJj8ujGdR258J4b//QrOHgznTRL/gR8cJtOZoKhxQ8jRpqC1p
z08Lr4slKpoxAVuoZquvUywdfwuOeXg72UA280bIFkz9icDeG849zNT4i2OozZDyKNJiKPpGq8It
AHWUxpxCdP03a3i/coud6w3Ls7CTkvP68EhKJ2g2vyU7TEHvWzzOtVCkGxd0l/QA3/a6WN14l6hX
LAyWPzfEvqyKNOgBPLNa0AVP6EZLSa4L/x1FQE3v+2UZx/yAYLyPUJhOI1akvUWqiJI0TyJeUsxt
BhMbEyhrOdK9N4hkuxP7YpxUKBDby+2MSF49cIgB86UPDuTStyILAYfkrbKyP9BiMjPX2NofJf0C
CWJpWC38eSaypHzHzZFW1rZmHmHkmlZ+XUSTl88wsH/jXWP5i5ZYKItLwtFPjMgaQxkpKWwgDuvn
m4BScN2ynTQkODP5zdNLQTQH6iINtJwNV8/4MimASTxKespUbgGS2qVJ6UqLClBsRFsIu/Zn8/YB
NWS6+5rNhHn1GTcMEKQPvSYRaOuF1iJGOw+1RSO4Xwdkh6nncsawT9WBUxMkHC+YRFI+xfK4hOGy
rqXxu+CVP7MtAWaL5t4+t0e1nHqYd4RL/z0xS2Ge7kKOavC/qNbTROtJgJXqLxvCxME/1WAPYSvp
DjYLy4qBQqKQSbBODel80ec0wK7MU4lujsCo3EGUkhf2ejDOjICrcYuaxJ45pJabUEwGPYvoNgfE
45OzX4aqFQzGrXkqRgMuaGB5k6sugG88Xm3yVZuWBT9zPgkI2LVoLaSeDa//r0XFvQJMya7RB5tZ
5UgLbJ7L9GgD2ef/u+LkRboaTheTCExyFnQHTKDF1QvqQTVFtr+rf6YVLEgaejFt6Hm17+Z5kPZc
3hQNDATCKJPjG1jnEiNmniJQqgcbVz08l7N3flQ2lJn/0ctLTbIN6R0ZkxakjaMZbdELbr+7ns4j
++8Z2IOt4AM8xeCl1kQZ7yMg8dHW9kUb3L+WPM+TU6rLwY11MQ3Qc3lb935mUg9HOC1/lPtGFyqZ
w74afGSAIl2Pgt0I5XNgtQrFMyJ2jESV/iHSlITK7y3KF9tzo/D3uy41yydL8P6ZBF3Bw0PIq9yd
nf6YpIZm8mMddSir3vixtmnyJ+CGfizcuujHcibQSth624zr2tHfbnqGRJyCj9r45/7LGCTAfg3W
5Hu/laoc1sNElECS7ZapINvc/V91C9qCM/DIzYOsW5Zm6GOVXrqju9YXzUKV/Hk+L01Wx+p6ASt1
pJ10wEa7lZJQAVXpTFJagffeurRymCaJpbuqRnOazWD3Coz2z5f2nQWFWEyMBr0XWVsa7Pz7QPxf
w19UFQSC66osaQryhtL+pO6Y4hFYdcxPmOG8M9/08aMVVKwMMYZgcJ+JLU/eFmZOMIJo+w3e9f0M
M5UYnAESf5evUPF9xBglCppoCqHdZTl7t1ywDrFUqJVoKInBviPqG9tSMWcsul/uNziCcX+Pc+Me
M4C0JbJSDW6AyXkTyf09knmctPctwmOTIMZErfRrZuuabyY758sRXFrqgqHiRC99rzmeAqpquNw9
OUVjhe+2MZXvrP/BxsMQjuaKPRbFJr3C3nWlOKPCXf4YgGUhprIG9ZCN0HrL2Zj3Hg7DVM8wMEOK
2HDLpRGAeF4GlGAQFugP8SukXGGJVnxFsA21WndPnkaA+wz9Z0+GjaQVG/GCm0u0nl13ejkgMLtE
xrSWENgHNFPxyx94+ypbONqQXs4PrwegKSe4//PyARyIinuVDIVZn5O6ORAUzRFwCxrAOOdKVyBY
6jqs3hQqLztunZoYJnVfwIJrj/O6avz4/uAkMJDujq+oLga8osQjL5kNh/qTLlLS+roFbGxhMRmU
SJT33btpT0I2y5ug0WRtjaDbB3IvB82BpxkB1wzlViIbWYr5+OM+sNEFmX/VJHzxbNEhvjUrpWHr
apP9zIvEv0Qwi2zzBwaNeyYRoAU5i9wPgKM2JndzeCM1Tm7HzUAULYX1fLBk3D4JbMf8f/8dcqm8
FIDxZNhE9TNtDGFPnkTfiZ4UPiHKMfO8rJYjbHYQNExkJq9Mz7wJvSth/4vHJOOVCN1iOr+TpCz6
YYLUTl+vcUoEKyjXQ9E9Ersfa1U71yXqrhGXlRGkwTv6kNX+BHDmy8RuKXNa1vQ5UCdRgcT2GS4Q
JaGIxeY2/wU8YEI1Wub8hICXbXbFCCS+1VSqbSS55zdOTgnru4oYEo+GkkV5z1jaqgtal5g54ULj
WnXRErSkxaCW2cVGbAjvk73cOINhLqXtcfJtFqpSNSW+NMKJ30NsksKUYkhDHhJU2cE01vH7Q3+U
adwo2xTZ3O95rFixhg1XcFWENJH2sI/kqZhYoe0Q7s642GiJVBprkjyf/IuMLviZmmYTq17hdVGT
7UmKDetq46/8fJA5tsZpzrKcEbqB2N6tcAXfppSwEieO39w4dTZmgavs9h9DU2YkVjFbREE/NbqF
IStJ8rnxJU6vS+AbXj4PgHcjO/5e3Gxsi1fhqvTxUV6DO6YO5H5H+DUNqNiBeIQv18QS5S4gfelb
/C5OCGMFnZKFiHcnIwyLL1TRSS1R/+fZZMq2FIIG4VxnvWZ4f6kbF9jBkiJWMh0IalzpZIGZu386
bhYPAmCSz5yoxMXV4z3vW2jS1VLsx615c/kcSF9Z0vIy94NJtV/N8OF7BdH+7cKSAZMp1iaU9wLR
Twfr8VHObb25ST9V8AVsZZl7bAeupVbpPUmBb4MX2qvxl32p1hvQ7gXRHUGiv4nGQasVy3lJVT8U
BoduOgGC3FvvVBDXSjbgFrlyUSspPE2vZ5nSFjWxF90AEq2PTsDIgSC8XOAI6B6W4/egaNWNEYXe
6ptQFKd40CCW7w/rd9eD15b+67I1LXNXIfxMuZlivTLSa1cvNGbS5R3ywV9NlY82o0xJArpr879t
dee4j/Ol+ySDVarfMAkXR0fBZUzInw+Tvc7VtoMugUyOfdW82N4/eNHMrH6SiTzzwcnF/E4TzH1r
6YKuNG+CY6K5sk2O79qCYS2MX1aYbjjoqB96Uq6Ph4eFiNR0439vAjYFSa5eiw7f/dHW5NV2QH1U
khTrOK+eevWGmDPOx7Bb0nh9BxSqsELh2L0tcct0B38ajtYZL7UYjkfuXOMgVNzln7xzNfXnIxpP
sEb6y5Fwm3ayZ+3sM1irX/nRPmiztqfpPEAsMcwKj1mhOjY5dG1Elgg0WZ0nn7ETjyoKtfPget1T
uppCLMQzOrTel76ghuslTwUWlqYDU0uLcX3XPZXctwfHqDRoFYot3vijOa/Q7AFURrZD+7BYujEy
QCKINlFvi45OxOwHDGApTLyxMrgWSJYJXsC2Ys9NbvdKeIqXhuj+s417oQFsbHhx2PhLU2TTf2uO
1N3nvX6YCDWCV6CNO1AsnhoItYwxDmW3JnIDp5qeGRWvpvLe9CTD97aw01j7UjvkdM3gZ7XAgidq
2pY3jfwmUUV1hd93ZEo1V3VRmGwxlj7R7TpIjyf5Uj/Gu3wehBEZFnblc4WvrpD5iP4YLMlZpBHW
u9fF/4Ayh6RfcJH8b9dHPzVjvgediyTOF3vIZiip8R9tfnEsn+rG/ftfpeYh6YHI6Qqk68Hp1cQj
1b9lX7r0RvnHfs/2hgkqrWrkKKciwEyw1WLFz89n/R5Q9wE3IsGL+i9cFZRaLwBoDaq3e6ed3VPa
N2Er9sX1cFlzl5GpOY1i9PaNyslkMHU4DlN7kRXbMP3MzK/6BFGYFIk/tLDg1mg+hyqbgIe9A7uJ
HNzNpUNO/CxH1NZ6kn+gfuVAR0Q32CsY1UkPLKITxszLNXHIkCaCI7PWjaYAKjw1XTg5/QblDtbi
BEsRW8kf4y/IL51n03YJ6m8rt96k5S1Iy4KTNJbfr6I87NqCV/gmatKxFuc2YBFYLbcGblSlMywX
kQOLjTWhbqeb0Csh9Fjy5JQY+xKgEsF2AlB9yCXVr04gfkmsJbm/hoKoQrbDObva+voIIv+TmJwt
v6Rw3i2reQ9bRrvzSDy+ZSkWPHdIYNhJNspUOE+8ROqOHxYfK61rRxD6NSjmR26C+LFiNOstOj82
D5D9xo6j8LE+t6Krxuom6kwZI4Ow4SDqa3S1K6vSdVABDuDxdv8gByRJUhmiXkU9ZievL8eCi08t
r/z96WO8ksNUBa91L1X+W8C73zjUqpA03fjhJpCYivLv6pxzDZzF5Li8meFKmRCYX30X+d2OSxhX
ij3Xq9PlvOemdAFY/Zgm7DugMSvL23KmajubxKfu/I58gKSltx2opSdbgG2X319w6hSicprzuldA
gABkluY5KH8sAL/5YnczlHe7yHNDNszKIHilO0ONrUnFzPrpU/SUo+nCtWTrcJN+of0PpvcdD9w7
v4Bj7xZLZRoeLKwsk+G611O5V3rm88AwyisOlt22VRMGNMYX5dXJ00sxZWjUPL0o9tut/ngI33TL
9UjjmZOiMXxpU+qPk1Ms8ycrx66yOeapvZz1di6DaK5saLoOu1mfzjOhEV8VY+Wa9FNwPrURmEL8
u9+R9hxHAt/FxV6VsyWWH7nQINqe4kBGwhcWm+8MptbiK62Q4XyB9Hs7JJgcPj7FPO7VpB0J8FG8
KCoyNkWiKDT2yXqjgrubOpnnGLfQGCe9EmkenCtElWrPbwwTN4jubga5aI8GssMeSjbBWP7IYP2j
7sfDwgMJN0CzZ3vdrSQ5eTCnJDDmYuLA8Mek3hc2TicuhsyvrPToIQuVfrBsDGC9+a3cpUIiNYBk
9W06p2oAtdQYQFPWoOIvP0IMhpPfrQFVKPGXCRTyoOmeKsZ84j03SYV0gd7dkSSdM1mohk10vhg2
vxVFiDH7olAUIXgPoFNBSH/1X4/sa+DWG9LVLByIQPylT+zxA+oiBB5WksXCJnUhCiICZUJpRDTY
GNg4p4S+i/4Uspxa+XPjtVhYZv3/SgNIeD2ZpnavwffeUSHqGJjd4evsF9Hi5VXupVWP1nUE5fZm
kQ6IIQ1BAJ3HO0kidCew3fc/RzMyG1seItyxTwcBfuQj/njKePnd48OuW8lchIvEaHOF+fsWbyeB
tdkpLwEguOkbkIVrDm6J+XSM8aod/YOygdiPvDCt+Om+E2K3rJxWnWLL+yjRhYO4jdB6N3jN+8xA
n71b0EfVLEzTpvWh0Ztc7m5n7vkIR0CejdBnCTCf6IeMUIWJwjAoTuvZronrq6ZWdbGRfVAkA/hn
F+yg4Ap6cwWhLioZYQDx1F/ESCKTdlGYCrIturfjOG+s+IJZ1toaIcdjBU+yovZgSb8neZsExDOR
htOvIy9T31Aku8Dnf9t1tSUDDJTMfVz9ScbWcln2cm/gByepH9QOUxHos/HDH/g2WkKuDPpuwdRm
m81g5w09tloo48MbdPxjiRcW9wo5/797kDUmGqr9f30GLQYlu+YvoRlRZCUwtInC4avZ/VhTt+L2
zzSEsLFUHAkGaMq72bhWTmYp1WOsoKYmDYi3oR3q2AHF8zhKrwKOLUv6/t1sSfAmIBJ8RZVVUcDI
qP+e9Qr+Qp4YXoLQoYpkLbR0JQb57UKceOlcXDiLrAfrJ7Kp4Ju/wnb18YdjarcDWcaraoVx0AD3
BgdJSdvrQNYUYU0O7fo8DSQClF+4xz5SgRn+wNRzM8A9gaw9h9kgv0tede83t3cTdNtkGoHWwcod
/aXZlHqaaHiYHcVlTj4/1MjL+MVEvXt0l+CTbCdMfjlcn4hYSNRiAnmIYNd1aPr5asphrSEmBorc
mQ6fLYeO+NYGLQl6tN7jotsVpmGy/hvptG9PT8eyUCdqCrdxR7jrvy1/m6ZGw5c/H6ljvy4SgyUE
77mfKdVAcC/59drMBimeMowVX97m6N8D3jokE+VCZhcdUTeCp78RPWHapNBmQxUENU+dXXnbW1/Y
GW0rFjcFTa2DkCnpgL6auOaQzWpL19PjbYMA3cEb9S10d2jzkU/CbnZamCuJgqjCyzDwm1pLII/R
zejH7LWQ1BNp2g/QQFPNRayQn8jKqs69zjO8c6FRZFbSi+03juYNh/sQSTBoVENJTeJpxVKETi76
UdqOm1a3r6akcYw5FIYR4XRbfLNA/Ze13MCUhC2Qlun9A4toywkOScLhaKzCWhS5DmpSvuD/modL
Udde9nrdtroOYHA7kPgSpSVrifuIfCgvwnLfF7I3b2VMCn/NzMoAfhgZFSMn1Z1NNexJTuibtWB7
Le0aaP0+v/1ed4lqZvIXZY0idSYILApW1sv5WDPzX4mE2BNPNwAyKP8LIIi1fXYWAoAHaBxmTx2z
DCABPJWQF/PnSr8e1BA+UFJ8t4gboaTEukNHSkQ/RiPxRJblBhCcg3GLY20h/Zys3zEOrnQp5OA8
SLkGUWK8njgwg8nHOMDcksyw3J2Qt5BxZhJYqDJW6nkjyIeEsxJ/nOIYY/A1z7fuAI8MuuK5Sb3O
H96kjl8/8JK/dKcNiRfP3Zi2va3i4inZB3d7w2TmvD7H5pkMsGbt8ZnBkJq6JhRnGWCBItYKYye7
iNPXl7A3CLhdw1dD0BqGp+apivxG4fCclPLuoGigs9AvlNb6F5KQ9hRHf0SWb5WtCzsNBQ496zIl
LmzCginBOOB8fSRCCS2K8ESI1Yon6T91naKfH2obD+93LKexd+pDH3tT/34euEfDJIENLFD6rgTq
ApSf1lcGbZRAcVETth9Fdtc9hXEYmSO0E3f9HyvPPFGXHH6Km6Dp0Vq2uQ+JHowsUhXNEAUQ5c9m
rkuED1bv7rTGWU8ntEM0PvSqZCBautYNiEuNOo2ZfsCvo5p76i69yeX3BeHmxn3KS+attPJQG14w
IjI0M3cXeRas+7KJdxuv+n+UlvOAs/8g2Ndw2LLXvUFraR1G9tl53lHJfYpzALs+Vztm7B7VtXbp
cOnaJiom+cwzotfBbSxzTT1iyHOAeD7CI7olLArjiDXIYlBh8PbljZdCCgb+oZJPvz9o4Rc/SIWk
NCeg6Nk1W5WyMJkWcx91j0GoB8TJq/V+z2mfmmGqUYSr2aDzfSOpxLY5Lg7OA+kVFmNW4VSHDmpE
B3nV8uwO5QwKl3Lc3QH3t5KvDVHvaNEuPSvubFnEPA651V3/yJsn2RcKriEGU9dY/ThGqasVt2qQ
CAYRCr3Op6RtMJbrUYlmsZ1+nxfZZcpn0zc/TzH8mN+ZJm6LH/CSb1AG3nEjQoo67q6T3KVVRTfO
2EPEM3qb5xWjdoshf37JoxEi873+NO+XIxbk+XIBpjTtvtOtc0SUKwTUBUOBZSyvjdSXAYRM/UVy
B5c/BgmV8dpKKogwQQPeFjsiE00CXNnQ1QW0LnvMr+ykLMEUWx6hSyzb2L9Ef2D3tFkJ48WTrmlQ
QtgQyKA1j+flpv4HtMfzpLMQ6mOvL/xNNYbPACcAxeeM0nDmlWu8PzkJ5KobcrwpBXdkA7kxrl9M
RyzBGtYTQbmvtsRseOz3gJ8XC/rvArQmu/EgQ35Rd6Sba+d5Z72sSdux8VTmR7A/qaZ46WOEwHwE
kqGfAp4XM3sMHGRZ1Hqxojk2AsfZWjaJI8oKO68YeG/DWmt3GH/GJDTlKItaVHyBEYagLWPiMbEO
uLNnIH2xiYC0MOvBg0vIl2dFBxZg3ARErQGViR2GobtINB2Ox0qeEsr3V25jJJO5krKrHLrIgwNU
hJ2xSAUjtOoaaat8HVVoaKkzJ9XP0eFzy8pJBuuTjc13alWs+5yfv91smaWwNp9GeMvOkxhG9YtW
APhuJZujlOIQoE4n2oEQwDZ5E3c7J39zDdpY3gZrHNyfhFVApYXJhhaQAhpzTpKPzOGEOHHJr0r/
nfZQznktDiyHnLIZF78lm5NsNhI7AGuTgbbV0NrPYSo9zwgnHqj8rfLIqf0A9MhEnqWIxkB4JRYi
rg436TCJ7vRTpBPuQLF4quHrkWv/nkuN7qXmzciEo3cOuD5gE9itx20ydi4q3WO+pvMiYnPfN0+A
776ft94UQHwsZozKkV/uSPMuSLgEqKGSrhqrrre8bcFCguodPSoK4d1CB7Hr/yzahQfkLB5Q4SNa
6Xyb3wUo1fiQfaFAgDZYmhE3LaQ588vdh047+0/nHQWtOhepbwuV0DRCCa+upgJDo6j0XIMhn9HA
EIrfK4gFB3HEIM8sa6O9/6b8nvWUUDODzBibQgQg8b8H4QwBOMuiDUB50WTbw4qWfaxtNk2FDq/F
A3zPjSE3951iWNuZOB6VNWjGiZ04lSSzzyvm3BwTL7f0Ci3iwGroLrYS4OB1weZvpM6f/HOYUkH6
BphCDp29cBHSfYpk3mgetHLE/xbyvIF6xQbf6G6nmz79iodmtsWC7nbUjkMnDYZqvOCMTGsHuEDu
QORKtOrQCsDcaJnNvhW/8e7IjT5XzL03NyW6LPSk1+vDe1jaz0ecSiR6d10S/cdvIgwnBYqQBDNz
vDnSB6e2fORUdYjmid5cB3ppK9atQ//lWlp8La0vlzUy+okvuuXjUmoUzpCgSL/t/MqhTHL/fuTI
7PIENaJ2F/fE30WDZf7YjRxx5KzC/VKZIU4yFL/sbmNJpuhCOwGAxtlS0qUNh0ihC/CtDnqnaLbM
RF2xNHIYqMTbfyBHfaYXbKrH/LbhfkNqIQmZTj0nCqBoS2E9rGloeVv2JohkQMlcF5OKD/VpVIdO
Y2/vAd8zXBRFcG7gVJORIM5IGg0L0TfFN/QCuQm/PnjY2DHsNNvvTuxx+XjGVM2SH9Iw1pPu0ldD
FBdF7Ci9HyR2luJcHVjJbYmENfiDXvCCtyGY2T8lhNw8o21aWrAGKdhAjGxVeA6e4NRstCT6CsY7
SF2Z1Yl0m+7drVvyjU5bYCr/rj2PtXxmvkNLcgfphGAp7Us1qMjpQEJ4kcuaKbXQg+LjjuH7R6eu
flZLyge66ThUPrRHeum9mRCqNGY9nbrsysQz9k4N4R71S+fXr8qU/74Xtzgmu0ZOcum3U+f0YWLK
dEkobO7X6yR8u6wpQ+c7+qJcQsv2vdqoqNLzQdrdEVsXAazNZUIgnlgQPmKHT0Ec9ZraV3A6ivpI
l1uI2h7Zz/YlYYseKeiD2G4xULkVPc2Lf5DCYpeGHdRYdTj/fP8hPMq0grx5ps2tmEC512soLLxA
o3UKUM7e/gu0PJO8sHzT2Ja7V/tbSZfT2htZaU4ICOlY9Dbxa+9h6vQWbZWpZEGMj03K/vFoyR6x
jZYtuUmYhVvUaD1HSJsJxwryks2AFGo3emdFExt5Jv+gREl11rffMz373fZju7RRi7ZpCR+92MKX
14uC5v/HdLspgLGKIzt63QvARBcayUsHJv0hB8kp6uAeeEWSe1ZXAAWLFqjngCnWeMZ5zYMYsXau
mR8h0kbFexzUBlsZjYzp7ar7Hsp2QWnFHJpt1c9Y4s50n31QHTUO0ijoe1PkgLFCYsn8mAvPSDdt
nqz2fCn/KIqxLpvoXLOF+VaDpYq1ouApl2xznHoMmhu6q1GmrMETpYk0nCfvp2Hjj4XDmVsOVP7c
9dcc5K+uMIIU263pB/kD0ENpqDWuAAOymiJGWIqOxDIuyszosw2orVIHB0cB4+lSNFGhoFN5n/d3
+0jWw7y6M7+XgVMNkXibzcI60oQB6dlcLQrRrKST4k8Ks+JeYzQWY5eor1d11TXdaXU3lJAE4Sd0
hqw5D+3tVeEWFIOlIhVyMAlOu+pQTJiho5YnciHuZT6mYOaR+IdT1Xofh5gtDLBty+vjU6pigdO1
FhCZ4s7315MzwGAf9dDbBDY08Nl82gRf1UVCaTS5Ijq9FQ6+4nSD8JfthHtCtF8BjO4OVVbiQIN5
vMsILUiGRsK7ZQK8SkQzBXNo55+Cv3IaFSkkEhtB51pjStJFrRNtAbiaQfbV1xSBP4XNmrSUyrWJ
ehXMpjHRwi3HdECKQp1usQIerwg8Jzik/JrealHPYWsEBU9KwfsMNRa+Nv4bg/TCIQ+0uWXOB2G6
eIto6IZJIM9eib5sZPH7gRWsvpZBsRwa7OThJFR9tz9GOXcxKjNdNNuHS1iKuJ8Bxg+wk1FoE8NF
TtOX5/eB2UF5GHNWJMpkLNUgdwYOD1gMtzMMshCvF/xVcMkMa7fceu8SaOfJ2QpYg8rTxtqe12/O
YP08MPB8902qao4kwAG6xURxkS5eTQMrSsv9RTRqZw73/CxOGKH7YEtdnVOZaEnmiigPVF96WvWN
7JxI+RxeSQJqia/kAEJ8suScoIDRW1zcpOUCZkchB+knAThbjeeGrG+ewbfE/1CN11ZHk/7mPI66
6yKsrB7fHrGBy80O2dhg7T/qPHGX0FG0/7rtmdS58dvYuLpJ5HusH/0bxw57LWmXfSpx5YzqzHMX
b6u53/7VNtu+Jd3PI3f0dOgPZbtNW5wSY2VfyjacaTAvD9WlZ6wBbpFaopeTdXqBDrSReOl5Xgvt
K3ek8GyzgNGVK2U04QtdtpKJiQ+83wNTaC9SmclmPoGY8ZlPLRr6XP1Pk6+Gw64fCkldgsn70C2X
cKl2LccoDDMBUmliqBXNNePV3G9xo14/dW/4sGPKcz/PudvZXe8SykoqoRpOrDSIw4Mhnl+kX2gG
nvEX+DFdF9ijDF3qfvWmEn33TmiSuqYYPw918Dk2OcMTvRlhPWbUB8ATRXo3IltOUAWRTXUd7nTj
mnkqcuw/N8+m+S/8xDYRP3MNq6f25y+dWMpLoLI4J4/XlrPALz1EdgEYv9/i18jR6t5SFRyhnL71
Rv+Q7wQ2RVgSBmaw/G4OXfF9gfZuPBrWsUXxWC1denE5xtur2g62Np+DxVyH23LMbyDrZ8PWVcxs
k+eo2qQEL7dzobkPpYAWLiDICIiRT83L958nVyW1jLnI+jziF3J9QUaRsQuG5Jma8ddDeDNDW335
SkzX6obeNwFzQCKtSCEXzwJwJoeh1pNg8rsqy03A39lAZC7ZhtEM0gbsM0YddKPPc3G/BZkspctv
ESVVxV+kcVeTiAyXw83ig78ai3XZan8XUPYp/4Ea//44uAGjldOMK24FOSiuKiK9b7ph48AS/SwH
JpXNMXl3ktnIlFuBgyMMAsmhnVhnrZCya/NRj2nw3YokpRyq7dr7nxIYpB/ff7OotgSBqZiSOwxt
WzdAjmxJKymkEApxob0dNtr2lLv6U4772X8bY5OU3+hU++NTJCYxmt9B+La1Kn3dVcNv4VymQv07
G3+cud27+7SN+mVdTkd7IuYMr8eOx//PCJEqDHzpMsY3LdxC0MAD0ISelYdyDglTOVa+R74ofwp7
m2s/Afz9+53pxF6OQzwBakSAQfoopCit1SZXboozph14/he3KssITW1nARGf25IY4sv0rEt1d1PY
rQQ8iRgDb1rN/ELdzmiBehmNTZtLDtGHBElVPlvuEV6Wj9bb+j3yPKpVBt8VuceG3Ghk/LbfWNNr
PfCNQUCKwHddCYX+R2/NIZKn3ooEajnQFZkY2u/bgh53dK2VtkCAIaygaxBh3KAeKvLRGoYudFHH
7ZvckGL+X4cGq0hoFKoghZPn+j5cjj4bikK2wcMl7C7zvJO6+8D16JiXgiObc+z3/cZwNy9B8eml
DtXQfcMMIspZIsY+eylphGdK5lMGAQQS7NEzhnqCURoNdJVMqX6H/1bLpMnY1fddedWkA4VyoOBH
Q+PWjYq8njjLhy2SmN7lpZQF0ahMfHaWg9eE//cron5GmCXMfAHROMxAHqTPiLaartgtYHSPmaBn
PserZbTOEhC+2qBdrTpW3pW+3mrIPEx2NLIEBbQdVpfSfihIZQ7ZpwleK8Rnj2ERNju/cWAJCaxA
Nz5ASF1JSxgHY3dp70J4o14BCy+x/a3ckQyRPFsKLN8O1f6SNm3qA5aSAtbPtQ8TSrdUk039OMvC
eDECAQ2Rux54iZlsT9XfTerYrO9DHRK7kR6w5LWCfpe0jDr1TMxde5b7zLkO2i/XGkeqt695+Q4a
G+7E9ygyT/5ViBlgroGyB6rCLW4mtg1e6P4F3BDTipg/1nKtZKoJBFRzIDCmmE+rxRo/XNSsN/FH
Ooq8f1WKCVLIm/6sxAxYcmJVGcQLSjmYBG+X11Zbf+QiIbkcdYfSukfW6uWfLvfinaZm5Jan4yjU
pqEbiu7RzDbfqzwkd82qiZGAz57Y+W1JxOCbUTf2T2mvpy0uOmoO9l9nw6w8EqwqMBxuaPkffn7O
XWkCSWHcjKYIhb9aPM7d0I7oisXuDvGNOwevV46vzJXFN+k+LYMdiYkulEL9wjl3gAqUkpfbowS4
sL1U1E1WjelbmYCNRiW27/9PXfl04wYKZfoqL/6tEKECe9Feybxiyu3PcCcWaISDj33x/jPV33I1
LckBZII8vV8sAxaEOWISohYnUr4HcjDsCqa6t6Fw42W4NSTDn52lU3vI00DQN86gK3KWJl2Aq6ce
kIjhH6pgTrk//gd7HpfAqbF8JaBCQjaYxtTRufRz1LKfTQ7Ixo5JG4uLZ5lauZIihKtpo76Titd1
CIF2/BgMRx4disfjOx1uHlhQOGNuyMLMSRdglUJFDcyu76P4PDiHoZUizaEARg3Kdr3vkLLyT3iM
lF2afNzHIg0PpcF0HgHFw8Pi7JFKBX1MLhgaYac9KNsnUILyj5HaZ1GNWB7+p1emUa6j/l+1JIkZ
eiP5DUz52qXHX0Fb0oRR7sYYknOLfwG9x8PoLEYyAr8lin2mwJA6WYkaguCHqxb3xs6C3YFwJMSv
88ZBGvCnAMesHkTInk7A1+TLgC6548NkZR6zXh074DFe6gqJTdEicue9pWzflDZlMLeMOQkozkIn
0NwrmP23cYMTaYG7z4yP9fTadhc4MB2ofiu3IIhlvEXUp5CneocHYIKc+LqAuKOXV9ZAH+25WdAQ
JkDbgY+Vt0QfTEz31tbzQLSuMwCdxTBu/2lZedSrEDzVRriEIO6xypq+z/ox1U0H5Yiy1LnFvJld
Nca2VSLjnjwMOxfnDCEjBFZgYSsHQJi2W1is700q/dH4IMpi9yFX7VPw1U/KKIFUUs/0WUHBcldu
EtEgf/X8bhsxFVcrc6exmeOPVDlMRXJ8vysvyjO6j4CF+vLJ91anqtmksOknPi1E9rKJCTb8pstf
RRGeHFV7FkZiH6XHEpVHwN2nryB0Ld9ykVPSw5tYeGkSY5Fb/xDjkF+NQ6zfAkAoJPtk/z6l2iMv
hgskk5HMHrDOMbxG1G6UmeLgR/e5rApWHg8zOnTK/Z51H8kUqFU2gx9BIKx1N8/RB6taqwF9PSKq
RCb/eM7rm/VovML9RRwDoHu+o0UBcVECeRGm0WSr0GMKNPm4RjprYinksjaxxh8mO9U17KCUaKb2
1jpz8D7s9Nm6bx2+iiDl59gcSMbJVI2tn/j2BWe4Xidt1Sw4mx2TA9dE39AgLoMspxqSK9DdZW32
UpAPCyBFuEJLswzjcITXzphzGNZoC5qz3S+ch3KuNnjA5uD9L719r3XBvfXf02vLcYCMrRXN6h57
lmo64Yh4ohSQiS+uH+jtE8LSekPF/SZYh1x5Y1d242x9YcMO0fB1TOZN1jtGTtnvLPGfGsnhxuO5
qFnTGLzDPXPfAza9W2XNU9agd8xkYkiS/ZJ+BTnkFOoTraSv4vIsLJt5U2tIkuUFdOZnSaSVvz3G
icmyJARt910JcmwUeZUUCNdX0HgaCaaZa2pJcX+xbiX7K3M6oX9MbwkEckjGuJB4/1c65GSz4coF
lvcDlojeaWYiiM1F6NhUahblWe56AOO1UFT1n1GZMhPJbl9jsXR3ewzQ9d5/Cl0jjNDCeAAGWjnk
Cn9LdHPerz515zPqk3qE5kdh2h3ivgKph9gr3jSGPqaVxGesbWWMr0hWp07CHsY8uWyChZhDoPf7
8LYSKmSGtX4uW1Swtm9OQk3RCUJE2+ayElESDszWsWktGwctHmeK+jDRpbBQWB6O9JmQ+a4obswy
WX3ttdkAGA7jvy7sBRfUJB3OLYnJczrcZkYTfAJ2LEgan7r8hsnTSVi335qnjvKCAIp9l6Atibd5
8R7hPK4bSXcgBjzT1lw1ZYjA+fvatnkMp8SNTyiSzYlPEV7w38dKUAqb3dHRbu52fgSQKaXQ86lm
8IJwRoFVW/kYPgn1AFpm+ecjfOTH6PUAoOs1R54hpyREQjiIYaespVY95/+Lpb3R+xb4aulMHMb/
GyP7elth+YjcM3ZCWTOVBnNtiL/utJdNuWLC09GdzeKAjKx7RaVxZEJCG6tufVmcsRHG9FeyeI4V
T9YwLeTyVql0LW3YWOfaELbPuaN07cOyqL8XncZFobQG9k5LoxAlFWTd/JuhCfzLARltWBg6forX
ztEHRfBBmgFGwu3b6Eir+Rfqx5z/jwcjxO0GwXE25tAWtOOv6HZudowm3/mq0lQQOObyqA5aOaH/
epafHKYJOKTbEdXddIxk2huviHnXzwoeXMTByWMRTfVgS7aXBnuktqB4r3k0+BkNrabSum8HUsDv
EA5rBXL0HmMEWhibF3Mnhl6X29OTa22c6QmcCihHCBunXCKQ7EfKQZk4XH9ef7qbMItYyqhQIxhM
cgm+V/XK2luZ7vLk1KBd0QxKsNXidoyHBK0p3UK6YXiCHebiWEP1/C5XdKyzRvEHkmknCcGi5KXo
9AyDmjptIhJhrPwVU9j7hcvZl2PdX6RLCdN7QEan1wwXEwEbWUNSOIeLYU7+zuX5xRJ/PwC5KiB5
Y+QLJxYWzy/2+4OZCBaePU+jdn1r/FQOK9uUMLbLbABLMdCFA59l7kngkSPJf82lTEk0ShgMrrD8
yL5HDKCdwQLDKXcLdMXmFMXCDMRyrKdqZYwyn/BpfP009kUvuQXEYTbrPL5acKwO4Hr7Km6akTxr
Wr9fPtjAZ7pCISwEZbpZAnP/o1+gMHBXSEYZy+J36X1bv1wKtXpTqftDZv+3+f8ive5+BenUXJBq
i5VsuqkvPBcmDrz7Q2G3yb/O1aae50ZPN1jemh0CR8oUqxJPfAM/2uKrjkPefy5bDN3rGRqsex4O
FuYw1LF3xvX065YX4drMszEMfviKfjDDvsKTqEI0yzD3A6LIsBH7YDKi0E6S33sBVEwm16BYjEVA
pZMKZBRnCtQIuKNXP1gjJyVf7+kKjYAJC5IgXJtBp5+UxycQzal5jYNuEN9ApitV37OZguaYDMaz
feAUigS9PEwP+OKp45lEzsCLU1lv4pN0td4bqRkK6o+YvDKhhCuOek6iG9F7bw50qTNWYk2Cl1pV
meIJLQFs5J842nPtQ7W108OoxqMVK1FOCzjQ8hW/F/dURVZm7IrulQcjGlLR3TuO/RyEUxSOMW/x
N0o1J4eQpx/qIKY25f8dN7G9dxpfz/7bDTVOVE30p2iufXtTsKOIuRKaAHR8wm0Xp0GaNOHKsgVX
7K3YuxOa+1Xe5LMtuEd3G9z23wQERzon1va62Lry6OIhjpX2fca4qWgvdoJSAuPxKCPMsVevLni0
rkiemPWcIE2lYKHm6vq63ZWDersDSSQLXmKWxYfL2FPAmDC3Od2AxvtyK1k8zl8N/I6sSXE7ZKzF
YVo6iGE7FycAG+4KIwvwL9V88bkGlA3VvI4LFeC7DLZmayrOZwDNpMfHF4cB8iwOavcbew2E4Jw7
I1KgK9he6qZ74AQfTp6JIwc89nt1J3hQDY9ey8lSepsDt5o3u82ckm2oNF/U0vylii0p2qKcMY34
w1NT2jmvuL0jSL5HvG5cAyn1LGXbwZBFM4g3e9mTNqbXmIzwA7dj72LpK3iuPYNsMzCLu5rVGb+k
EAobpd5PwHGk/kVnU8Vzde12jo0Y72JPOuBifrhOtjdBs29jXWekhh9pY4A1vnOVE3zLVQfUPp+q
Ggm+PZmnxCCym4WwafAaBmblkXbDgzoPh9iiHg9aWRVNbdM1zpOo+AWX6/kU2zzBEerjVNhDEaN3
4wJA7kOhxSjfbr7/DxdhEsgRYtMweSOJbqxLAG+tRz0gVg7Y6z94hwibgxFRyboXRHE6C+QXVTZB
TFBIrBa1bQ6JUv91hOLdU/DNDl1Xckhgs191McAv/hGEA+JVdvUF91Pdclto72TRrmg1XaGw7KLb
0Hu8EusHsDLWSyKiDka5zA7iV8GDNESKIu0nrqkozxZdKvS02CXlNBbtkAD2sYVhIELJuoYqGfzo
bo9IGVLuKgZt60ZCxd41yIqSbcOwnluxrEj1CxZ5J4L9CVzRk/YNp6xbrNYM/GZoJ3fIkaseionB
MDDTMZ4wo5vs1bZm1CSAEHra8PAQcKHF288EU43CmHiQqAFJ2JCzznFLEm1+BVJ+6+eK6zXA/kbT
qIMDJxbfdnWWIOKkoJMlMLGCRyOXCi/BXQCxQuoNR/pc+qUntArA85zMvRR9BF1ut596CO1LnYvj
D2VMoK058/dpEEMr5FkeHcaP2tlo1CEzdjtv1xPdQp28t4/7QpxZ59+yuxaItth8YqZyJPF1kYKa
9d8ukeTtp/qusxRLiJdCxz9iNZmfPzB1HA/i6VvsxcJJtVQs7aopkVzRkmBBds2R1QeRE6gdvtLS
6jtgaRsc2RBjxM20FweQjTyCZZcmmbn9vmxyCdclS+WdYzKOldYw4x6+ksHu7oq/RYq+lRuPMSHI
l+UuPP/LR4vIXRy19E0VHxWOh4kS+EyHLA7BuVfjKrV/B7GJ3KKPl7sw58KL1rDpR180NrjkOFtx
LsJDVrvBxP2QzPs1faREbKi4XXboD4A5tepgq5R4D11Qim46ogWTcYfldl3AnyTBdvcBgfz++0rh
saAsA9MrAicvNLqjjMm0nJDqjcNwthfrnGP71VMI+eBl9oFIadCuMtdaKSbdfZx3pcjzGyxoyANZ
rzDv34Z70tVpMmnbEZ6up/JqkU4N6qAipgZGyi+T0ee9+wM1aSt3+UoADLpjNDD5BH8cJilMOOkM
d96k15lsnJtkOtVzRGDvLjeBLDmP3lDU/7Zf4MiEVCt9pBXi0e/OK96mCturD/n9AclkrpvssFNn
GDju27ENXOhZtiYKsMyfnx/HYRItV2V5BTyzdxElYHQs/3cX8zxJpBWKkxRjLz1TQAIT+kqo2C+2
Rh3GYZ1Uy7KkMhlnLC31S9x3xo8fH2wr+VmUxjq7zCueqSkOCobyzMr7b5qRRZTQYC5lSc0o8my0
hOjy05qQtDI+xEN/4H7VEvhTHYSX7sgco3Dt16TictLl/ZlTY/axlkqPZ2zrY4BdouJwHpMiBCkm
42bz302r6i/2oDSpQSUGB18ntg84O0togMc8zPzaAPQ5uiWUfzJPvmdJXWLMius7X2OxigKSpPMD
zJlE26CMU2ywucGx3309Gfpx0JOZiqD40JwTHYWf2spLI4jknNSflamJAfDHtzx90+rA4hz24VpK
yH3kK+v7xmjDKF3SbH6Bgz/xYX+34q8eVq63ccLGqxayWh2CCdf/200zNITw4K1OHkdGaTO+tdnv
a+O0yF9261ScIJle6R0e3+lM645Fy8mlB7HZNQEx6pm8ChqQ/V1f2RZdIycdCgCpNkW/2kDNwLHn
kwJGeB+J0NgIVQHgAJPg2u1+8bwvJlYra6yCjoQiz+C7rdpKwShgnHLODfy/MhjA750Nl+P3MLn5
ql8skk7C9fTtukKi4Z9Ce58RYgUbtZ+4PgKxmxp03VtaXYK1OBrb6nkK0cI62DDwuDcjAuWFBjPu
lAvT7d0xcfyFpAmgRhtmLORJBs6fszsajHgfaP71zJS5yn6GU8noVfONeKp3k5cKx/6yfOkzj1in
uMdsp5uATsHp9CfwTjzWcBdAAbXfw+J1v+Ja94c8XfQvsphlPZDKMYn+3RGTBGyx/QDk7eQc2g1M
QBCwuvoq5CQtDcKJqmCbsEfQZF9z/AYRtpy2/gRoGmp+Y9qNOVeXI7hoGtftbt+ktwSlr3qRBbzU
nKI5jiSGkiuRYILHMeplNgFGN5MgRREM3kYfiDyIQbbBa+whTtOmkq2FjE4LebQYYw4AThu5oGzX
QLrxEEZd9/md/eE6Mre18y0uQl26DvqUXzAAoGrK39/mRXdIU62vF/VqEpc7uMuHQrVTDpVCy2bO
hZND2yGeq2bJFQL4ia5zvCGk6NPfYe2ce3hs/0v1ipufL+3t6+iQ1Or03fwPVF2/lNX/qM1zMtc8
kBXMrMT9pv1TEMYkikHmzk/oK0NFKKkKB9RUvmRpQysPYYre3IpG6erlCzthwM5O5rK+5uZ3M2oU
v38MXRegachr1AgTMfn3iqGA3W7SiL3nWVy3yD3GtRqlWafMz2Ta8X6rHEeXUqIPoHLPXiBI5N1r
qV55pbir+zffvrVrM3jO8klS7jibY8STRjFA6on0R3zhuKHoSzR454xDMsoFCE2cNIDN8HKBKvdn
WYJZwejhgpIkThI6rUJ+zF5zALrqgJIGIqKAtFteQ44f9Cv6TEMxQbGT/y1790ZIJ+jzJoD6Y29U
jzwBWJm3FIwO2DamhqNNTPXY9lJaaM0vuZc1XDkRUkNY5TBxv0XOmv5Dkzyg+Ti2xO7wIyon2hxD
TBVX/kSBy6d5SqYESQUoFEDZQb70R+PcyuVzBwCb+FbeRQtm38zU9TltkKiD0RxSQudYN3caIYgi
/HVNTCqZKEzYyylnzn0NWlcP848WoAS7rmrGmBvy/kFaNV30E8bja4c4G641DfSrQkX2yRXVXfgo
hGDbIcYFqTlb/yEqDzaRHLt6+TcwXvd9LXnmKx83rMk6Izw0j/slTJ8fdpgKe+UBAUhF99Yx87C4
K2Th6rCz8Ni7jL6hWOQMtzHqqPDQq13Qyu1Jt2rqfVagRC12eqMgU5JMfsJO1ifpEr6CK/yvbxI1
apxso/rjUj6izGLBP64krs6BdkvskNhTQlCrRh1y9tWZ7crT/hVk3zCYr00aqYcTLrby1ebcZoc4
lUCt/1HncXjhfG4T7TARCba75puvoSYCn1cByFSfkmrmrNW7wm/z3NzpYuHsT+LJZ+D4VJzyLw5o
WknaQ7bBEdzC3kusF79JY93sOxwHeFuKQR93ZmNHz2zPAYeahSXlFuZfhREqz1+Zsg0m3aQ7A0kb
goA2irRCYr3TnCe0V4YDtta//52/zwt9zW4KgtYp9IDZrWcTtMzKchTCzNT3L9VCvegELt9C4ltb
Nwh9yqoJaejG/SNg95NfZiJyB74Q8XqRMlykNm6NBBGdFuYoLvy0hHEqC0DwBd3cwEVVkTn9bpD7
a9D2J+IZhJgBZ0KWmxYentYsl8sgJ7XRo4lnZu1Kx9C5GV05OqtyIMMeTkI5kyvhxczLWjQVHZIi
rAQkTF8SrJIvhlgcbjSkElutnPHy4zSxC0gMtYJw6B/MKMb7WEnBWfNSggIMqWNoauwoBmdL0Bcp
FuaZ3EEsa1tdAZKbaxV3vhthzkRruom4HlQhq1HiQWiXffPgNsfM3UYpdXjuGfQuxo2GTW2ZKPwM
83LWTkK+LUaA4d2g5qKfuuzv3qug9ndxNj7a+ynMnbsvW1gtVlhvCDAtP3/1mEpFmDiWeC3TqFeT
jirWEIp9UHKJgi4Wi+6VVsCXiHySpNy7w+0tlsQOKPuga0Z2TRwSFPCG0ugYZ+RgOR/mjJI+KBbx
nPThtm8cWlikldIqd87LljMuSBhUo4dShZVrZAPEbFQrtppHxeul2e4LYZsev5tPtFN2H91fDdtr
gjqgxxeKFSOwotSOQw49JXDHJAzudfX+9O8j7S0czYKy42wEy1pfh4e6cKDY0FuAooXar43aJNmo
KawrD/DsQqdP9lXgU2Yo+qf5NL9Py8FyTFBrxQTJmBr2layja23WotfNXW7wIWUfJzIAYXIjFzPO
EizQl6e6E2yVTDmzepnwZhlCEGJfOvbNHOKtfLXuuTA0yd54i/RcjpBIRGVqa3rK3rmoJCiPjer8
ZimlWV1170EaEUDNem0BWWs0mGxL4tgOZ2Gmbv4kYShD/BATX7PAmDyoZtjw1mD508p0lbOS01EJ
O6wC8pepY0VHJ/WHpBNoPxl6Am9QNj5UwxTMzEg19X8NEurlxYfG7wCv5PYPpZRCrwbxGPzxE8II
YyI1AEWU8BX9I01/rZkd7YZtiEX1MjwoQnqakXwfjW4NTPwi1U70eUQS9j5X3Vk3kOq9+jFevLmz
WN5qYUPvtfDpCWMOIDneFkqjKkLVILxzJsYhZtwdnWsPuYE9fQMwl6EZmqN859HSEdspSgxK6wtB
mUnz92Hph+TwjADMXbBYHBiKkEq0TAFSKE+rpN4XVE7iQhSW+qZ/miJpPzeGUPZNAA095muy1Ays
EsprSuSdCfENC8NZJanHGHkLMvkxQ/ypeU6QxV5xCU+Qr/vW6OWiPLgxcl2+NKFmy56tCKKcxvYE
OaApErOx89qE+bqCRie6yHLSz57YHR4Ex4rW2XPyKxllpOFAPCkU5i6CTUZ2mxQVgxHbTrPNo769
v04VwqOSWmoaQtT6DmuOGuSWBdV56QZFiibcLyGC5V+Bn5Ew1GJO5pA+U8jF3NX9VFsO4uLRpE29
O6emPYdi4YxqqZhSfrZYLI2NOfHjsnSlAVNciWJk382m2R3RzEulfbMUiiCM5RvhPL+LX2iplad9
5xDvKw5RyGvkrgZCYGiA9JhFicwHwvl7AKLB4kfIc8BBmv3BkDj6MIiTuqEy7kcbvBqDEO6PddBV
KcbXEn+gFLNzPcjIl5x8RJApi/TzSOn/78jkkckYZWYroz0GYJB7Cog/TKpf6sRrgH6jU8MG8RNp
x22Wedbzd4CCG4m9rhOGcamhNJfKJtel2r/jE50OJjJ2bANaPpw3LvelTEVhHW5DY8KwlNfJHExH
Qm+fESd+2yOuajOf/Z1If07sejlSc07/9NrbLlQHyWsUHpW8cQHVsuxlEpSrtzJ8JsSNTYXAm6PU
eKfzubMVD2G3teRH9m1Yf/PEob8cciOI+1Is4eWLa0S0Geg5d/XY0v5u/ZyoNVzuXkROhj5oZw8P
lM6nyWpK5Thi/I/ux6/kJjIPI21FBxaWD51YjLwimw7X6OVdK9ws0kjoySwFBEuuevXauI5xv3jh
UHY8se4X1tggy1ZhZU3IrMGWvJDXeWhSsS0wqA3blVTTLEpvRGBPLiPgBrpmrC5bSifbaAR9hEQr
KA3ePutZKCCrqvPHEeqCM/bsXzi+SMowJvl6pmG7uA+Ef4xtdQavp+MGBMuR7RAc/8nA4sCNgAmO
nT5NBfQ5tXEfKttH4xVdq3jjvjBhVzP8jsnI6zsRn2be1p9tw2XVg+OcS+saRcN8qfaAazucWccs
PJPHwo2hN/57UIMdiBLsYSY3E5qGtuWv9qReq6AbrfGxIblZWnThgl5jTH01TKd4ExjIonRL749s
uDPE9ZJ1ISK4MhCEI+3h4MY7LvETlSVR/Knd+PTHSN29E21dXSzOGINkD4IjcoUMEsXwK9qY6qYG
1ZcKkaIwjYa0UAhq6DRcVV2rMRVSzarZ6IctN4zjwn9CYTGbt5h+CMak3oD+JHQU9lidE6uXer3h
n1vztlzQyg6Fh40cRm6gbSlNO/Ouy3HQctak+j5uKbPrD1KMGgoqDRNIIk4LOrQMjUIdGbsgM7ud
0DJd5jvn79PrqgDRwN6Ougte1XfBq+ZsSSpPX/63jp4Z3hHazltLR5fkDNhuJDwg6Hac0Mqhg6we
LEo0l0nVYmDfQJfzzA31/NFj4wgfN1G64gDEsUrWpcgfudol6c5puWNuzdZOZOpl+eEyi0Xh2cOJ
t0YICiRYhcBPZ2q1cl/TeJteXrQ1PCRWQ+418F2Msby5nndfs8w9A4GLpXKPM+j9AT8sS5cP/6/y
nuM+NjbOaSraFHA5qJfY0Wcp43WOs7Aew0GbXhmgHKDc9hoYDIV2coYBeqH9gOZ4FUOwo56b/AFL
kJI/BoP39KUFH86mkJWhaujgn93o85bIBdsdS99RYeWpHaQTGqveUYxGNycts+zMIfS81UUAiNIb
f+ip8qDS+f/drC3tjmlu5HsyXDdwBNOYLknZgLfpKQnu+qpNqpnM9cA+BHKAd8bcTsa/wcpDhGZH
VYAzOMkKojY1Ni8THR0fdfuKXQXtLQM2XenyK+0YU4+FJDIzcjE6S7UpHhGjc8q2rwHnRzeGVVMk
I75eUePHaqrfUMmjQD/5z3NgJHjnbcPwD8Qra1fGy/3JOPMfrsmfk8V7lSSsymBhnoYx4tZKLFSY
ilSxd8ni4im57cZ1Qwjam4+z8YzOlsynBxR/4WZWOTrrnpc5wc2p0dywdvLVwqx0X6f9nXAZF5oc
Q02/9wVGLweIwMY8Pkci74R4Njtrq4caO7qVklVKH0fAtp1FIIgg5jbc29vwmbfwhyX3HClmD/vg
xYwdGQecwFdy3YucT4hgZvjLLYCE4jxht4C4YSIsjiHBI+r40CwwkelwGn72lf09nVjXfu+eB3QJ
ENRWVa+MoFU7urQrc2E3+N7+jfqSo8cohiS+6JVbrCtjzey6NmeNnzaiiDR00u5FfbaVzos5BluE
9ATKAiY/Gdga/UI6mlmiS/tYvs0rekfdMPNk5FMdw6PkFJ8kmS6f3Y9ro2OZ/CnBPTQDZQoOZ9A1
QgQU88CCRiBwP6zY4etspn8BpnRFLSyhnQTEo0yTUmngvxOm8JlU88dwcH8WnsN2UB2Ith++CzbY
/f3XUNi2NgnU/mDPSQjRPcWnMDMQMhW6cDhfnE5aPj0R1XQOkifS2lehjW84oBoeXgTiizIdXyW/
cYaYhBN7unde68LHpWxtrasKGNSSmdL19J1WYsTcYHhiVd1xxdtsNOJraR8HZPMgvMDkNjDpUyOy
QMCdal0XL56KM3V/3I3kItH5g+lIkCTKsim8K91XVDW/Rx92WlqD1Hm4i4C/C2sWIRcWB+s55iZr
Rkyoq2ptOwJeg7DvNaLsYdc1ks6ffRAD0Y6FDERFOmjwiPixbMrLtnAjki4CMTNPl6vj68P43PzS
m3FBEqypnl4POlX2v8R3H17+KxWxXcI+jTmScZ8VFpfY9VuoT2ym34kRqxbllqdoTIWFJ4f/7eEx
b5frb28C003w8xXGbsJFiJxUMvo0VSpARtDT2yR86I2xT6w5ISqYTWhYKebQhjv7ag3Oj8H60FO7
GIjcr3P+3EFZyodp7LfRsBLrRnu4B7cKWXo/PEkF6Sf7WtNpThazYXw+icaQWi7vcGhgEVtHH+4D
m8Db7mzAAJDQtGW4ui3dMIZ64Vff/fVuWmWbB+2MyyO3o6mkIqKo3p/UvaQvq25CZ8scm5OunQD8
DVQSuSZpSGEKz1uEAIMJWRP6PD8uZYEMs3TU+EP5SdjtOzfzhyKMSIkssYiFFuH1OXPD5ZgYbGS1
EY5PAqHVnbYZH+PC5O1Cm1U+roKCap77vRMAXCezyGAdCRmIRLASePLDcAqsuUy0wzqgfTEsOmqx
5gY1ZTiuKvjWYT2hr4/ZXVxhK2zRvDfqpW4nqkLFZwYO98qCzUCdoI9cjrgstKMvdPvDmwHD3hBG
WBVY8xohM+PeBZw/5Wzd4i5F9CxN6sfmtC8ChmI95RHBDToggqCAgkH4Xy8IsQ2ajIizr6WWvEbr
YA7TLlDXn45CtOXjKzK6+na53oAPf3UymNDkNQmo6e8hWIRV9a70CRilqK9HQRYHB9HTWAWogJHw
VFkBMzEx6p/+3wgbmM0Bu0/ysVETX6fuIi+YMJssrwqNKO8CCsw6rBWcxH8vP0kaDQ+m1c1z2LUf
pgavyxoU8f6FCofLun12sYvnVlgWHiHr5Qnaq+moWgshfanPB9URa+D05iSIGs93tXAEQW/VcJAm
EDUtLHQgfF2JBwoy4k680TvvZKiTSO8LaO5dfvi3ZFVV6laA65udlON541dDFTyp9v/pVz8JgrmA
BVs4OBTCWCmw5THNy32MIElZcacIeo3YGYE9LCdZjNRzWMeeVYcRypI9CQenai5cp0Dlexd/H/I3
NjrB6+zwMSB4CmRD7vPdZcWB/jPmYff7gjivCU/L0EfW+9V8yY+sZw7rl8QQ6UiCCZP7TwshvnvS
a42CeYLBKvqBouxBJkisphtDHBIHb6ZzJyqUgKyegXQ9B71ZS8BH9uT1sSM3VD8mEbv6hvonBKKm
Q/UbKlh6IeHNZ3vZFpohO+ZEcPKqUpBPiPTrD9F4E6hec1q2YzCSxNkRfTnGmsrCQ35IsRbkfvML
p/o7NpUVx9pkzgXgb8Jsd2ZBq2GtojvrOCuAq2YUam6xhjV1q2+tWcKE/fzKXgNUWOQXfiZy8Kfl
+S+e6yPPfpCnPbihPS9Y6rnKWoyJ/0OWkOpBq8Y8GnDOSWztrh7sT9A0nYizIeTTFaaG/ZcBi7gP
ee6RctN5mB1UxvNsM5CLBA9rvkPPijmVUAHFBasKea4NlcmwKSKFsC0bcVcr05cnG+1sPsQUyb2+
sooo2CBp5XYNSvzC4PGygxrMF1Ef5ESHbmWRJnB0YkeNoWQEsk2I4aSikCh1URh3pVvAzoBavNfE
o2lWtj9N5VoEy2bUkwsLAL3F2+HRTL7GseDyYja5TW3cS/uXMIur4v1xUCF6T7bRPOzoa/cuW2ol
jUFDK3mUsMAnvbObJJ84QL8+nKr10/vYj+KOwsKeSoDPMWIn5TGs6EU2E58o5AKSpYyhigsdNU0o
fe2YNNNHg/Mg1W3tpOzJW9UtvtL7ZbMA3u8oewKjtoF9MyV9tQNXWvNjcKvx0yBFP8Dr7epi4awR
u7hx4QAj8x03psBkp96raBe04zDJIcTBOFaWKHC9yQheo/R/N8Hnwq39wT/n0rD0V6CK0VmM3tgT
a4DU5/8r9C8bfQEg21i1g1LGofKeN5EqfB/xcj/O1sUg2rO3AhLjeIiejPhdZeRLHeHB5IlPf7o5
0OJj1Rxs/fZYl12SACHNa5fslDYnqwaFP5z8CxQyL7PpVBJ9chAZTS1l6zJIPUyT0cPFugWtS7vL
XVtjA7JNwZOOEFLm
`protect end_protected
