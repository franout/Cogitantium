// Register NVDLA_SDP_RDMA_S_STATUS_0
#define NVDLA_SDP_RDMA_S_STATUS_0					32'h8000
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_SDP_RDMA_S_POINTER_0
#define NVDLA_SDP_RDMA_S_POINTER_0					32'h8004
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_SDP_RDMA_D_OP_ENABLE_0
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0					32'h8008
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0					32'h800c
#define NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0_WIDTH_RANGE			12:0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0_WIDTH_SIZE				13


// Register NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0					32'h8010
#define NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0_HEIGHT_RANGE			12:0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0_HEIGHT_SIZE				13


// Register NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0					32'h8014
#define NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0_CHANNEL_RANGE			12:0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0_CHANNEL_SIZE				13


// Register NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0					32'h8018
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0					32'h801c
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0					32'h8020
#define NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0					32'h8024
#define NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BRDMA_CFG_0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0					32'h8028
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_NO			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_YES			1'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_RANGE			2:1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_SIZE				2
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_MUL			2'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_ALU			2'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_BOTH			2'h2
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_RANGE			3:3
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_ONE_BYTE			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_TWO_BYTE			1'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_RANGE			4:4
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_PER_KERNEL			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_PER_ELEMENT			1'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_RANGE			5:5
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0					32'h802c
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0_BS_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0_BS_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0					32'h8030
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0_BS_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0_BS_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0					32'h8034
#define NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0_BS_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0_BS_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0					32'h8038
#define NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0_BS_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0_BS_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0
#define NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0					32'h803c
#define NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0_BS_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0_BS_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_NRDMA_CFG_0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0					32'h8040
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_NO			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_YES			1'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_RANGE			2:1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_SIZE				2
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_MUL			2'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_ALU			2'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_BOTH			2'h2
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_RANGE			3:3
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_ONE_BYTE			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_TWO_BYTE			1'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_RANGE			4:4
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_PER_KERNEL			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_PER_ELEMENT			1'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_RANGE			5:5
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0					32'h8044
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0_BN_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0_BN_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0					32'h8048
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0_BN_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0_BN_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0					32'h804c
#define NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0_BN_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0_BN_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0					32'h8050
#define NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0_BN_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0_BN_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0
#define NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0					32'h8054
#define NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0_BN_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0_BN_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_ERDMA_CFG_0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0					32'h8058
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_NO			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_YES			1'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_RANGE			2:1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_SIZE				2
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_MUL			2'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_ALU			2'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_BOTH			2'h2
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_RANGE			3:3
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_ONE_BYTE			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_TWO_BYTE			1'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_RANGE			4:4
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_PER_KERNEL			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_PER_ELEMENT			1'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_RANGE			5:5
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0					32'h805c
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0_EW_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0_EW_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0					32'h8060
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0_EW_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0_EW_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0					32'h8064
#define NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0_EW_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0_EW_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0					32'h8068
#define NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0_EW_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0_EW_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0
#define NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0					32'h806c
#define NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0_EW_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0_EW_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0					32'h8070
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_OFF			1'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_ON			1'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_RANGE			1:1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_SIZE				1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_OFF			1'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_ON			1'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_RANGE			3:2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_FP16			2'h2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_RANGE			5:4
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_RANGE			7:6
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_SIZE				2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_INT8			2'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_INT16			2'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_FP16			2'h2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_RANGE			12:8
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_SIZE				5


// Register NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0					32'h8074
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0
#define NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0					32'h8078
#define NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0
#define NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0					32'h807c
#define NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_ENABLE_0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0					32'h8080
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_RANGE			0:0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_SIZE				1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_NO			1'h0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_YES			1'h1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_RANGE			1:1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_SIZE				1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_NO			1'h0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_YES			1'h1


// Register NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0					32'h8084
#define NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0_MRDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0_MRDMA_STALL_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0					32'h8088
#define NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0_BRDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0_BRDMA_STALL_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0					32'h808c
#define NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0_NRDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0_NRDMA_STALL_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0					32'h8090
#define NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0_ERDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0_ERDMA_STALL_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_SDP_RDMA	32'h8000
