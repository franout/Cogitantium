`ifndef __DSP_USAGE_VH
`define __DSP_USAGE_VH

/**************************************************************
	dsp usage for generation algorithm of mac units 
		in the mxu core 
	NOTE: board and tool dependent and previously checked! 
**************************************************************/




`endif 