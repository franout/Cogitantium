//==================================================================================================
//  Filename      : tb_dtpu_hiear.v
//  Created On    : 2020-05-09 23:47:05
//  Last Modified : 2020-05-17 12:58:32
//  Revision      : 
//  Author        : Angione Francesco
//  Company       : Chalmers University of Technology, Sweden - Politecnico di Torino, Italy
//  Email         : francescoangione8@gmail.com angione@student.chalmers.se s262620@studenti.polito.it  
//
//  Description   : testbench in sv for testing also the axi protocol outcome
//
//
//==================================================================================================

`timescale 1ns / 1ps



module tb_dtpu_hiear ();



endmodule