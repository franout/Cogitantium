`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HFXM4QpzOzpK/fVpfk62dyKPaY+M2q73y7kMST3Op30ot5NvOq0U6FCld24uN3mmdEOCB27hKTuZ
pvj74DeWqw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hxkDFNzsdQeNRsfOnWUTHNFz19Fie2E9Ww6bJtv5S8Vni8wJTCDEWn/VYPY5k60HVYU07IHi/s/w
GjOwEwynUdlKjmKERxlFZ0a2Yjq3JWwUWc12cFxPSFvHMP9QfWTysUCHYJ+8/RIfZyEk46bmujim
y/VHufEI5ZXO4q4Gyqk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ONAndknOfQIk+swhizfY1gL0lm7OhwKPDqzujw7z99+5JAeSmYF0iR1qz5EwF7eMf5o+eBBTlTY2
NjtC+ofhlJj3YLY8Lkd9hce1iIgbgxAHpNhAV4hxZNKKlcUJL0kmwJ2sBl2MaOhu9WOIXP/gyXyN
CcPlRENgwlBbU1+C+1iGMMh/9KMne0a6VUr1gNN9QtCYdyQPFjA4dIq2FMmTQiiWUgkSyYCsCyDb
DVO79Ar9lZt0fdkJ6i5QqmM36MBOVzBWCBvI2axI5+7vCpi1BqmzIplWl5EiE4AsRQfOI2TBfUtP
yEOrYnZyYIKPzWZQlhtcVDoxbaFCeUvUpCviLA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TaVTZb7cDJPqyMly4kBtJvAOCbKPx/eKng+0R1rQMo2o8SuEfVFk/6j76zwZHlOWuJpku6UpfFwE
plsdbFjrNL1PGJMg4nWHYsQ6cpSFGCrzsH8ZoOcnNJ/VlLa73SPXwczEtdZv9OKf3HFgn9MY4CrQ
2EawARLqvq3NHrhdYvp5AacISwij7ZM2qAX68EevyoorF63lRK9KOcAGhxo76mjzzoSFtfSjmWx0
JTymJkTP942KbSf5k0lqAkiaLOdR7mQvwPS0A2G0q8VAgtqOsBEluF/6E8KYxtj+LL9wx3GGpsBf
QLjO+0YsgDaQXX9OmrJm8KCaDRkoDHcwWQIAhg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jM7OeRTJZ5wFD3zH4AZkUK7T+3O5+GGAiKbBdDc7gC2sdtjbLkypvsOJC7Uh9dgB1Wdz8Gav74SF
K0wImUoQx9TOwcwEZjzl61xYSVKhdG13ztjZ8/cWPFwmBpB2uXVcFQ2gClKmWpg0qtU9W5ChP0KM
r2p9sLxxsNlP8BNDQLwU1SF98kYKf5AYdncwY86TqtAes+iWDkfIwS1+XGps/Yx0i3oh3FMEbNph
RklthnIT0OsXxkuBWmFrHLjiJeEcVHJJPKi3uVXa5Jt9ePPqy5sJzhmC/XCqNXSinsA0SATkrtbI
zz/momgxCWatRufAGv/asXlnlfymv2nMCYTe6A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NcdUkKdbmEUn+isQuriWZl51sQWsKh1eUDZxUe6WX9WqSm+N/500JA4WaaBP0pn3NXrK7n7uDwmj
4Djz2LpdFbP0Ymu7AzHFHf0IWC04c1QzeMK0yoU/mqVN4ns9sRIO4XANEka5JEiWkWlEasGDu9CS
/fpSluQMMHBSDGFNwnQ=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PwjOwv5uT1gLFZv4b6gD9Wm9pGXWuC0z1+Q/cLO3k0wfMfEeMgqGcX2tv/sky4agZcCf67zXdL5F
GWKwiANORqW8Y2DRguQ0Rr7qMb/sYqzlgoL3bpKQrJqAnNpP4UkUcLJoP1VW0MZiCg6waiV6ZF74
FWYgMBG+F1nsIpwvonUgsrZSP5k6Qtsl2nRB76q3WgaErOtvbTjA5zBTZW6cnlzrVEZYwHTlkg1D
9yVDXO3GLl9pvSCZxZ0iZx//96llr6FVgBj2TyO9q8hSStpn5HYqbqW5wc+JckdlJSDIu0p3GOQv
QmkXkkyQUZZyLCv64ddhIyW/PlMrl8y+9JZdxQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DuKwWtfTc2231DZXJ7uNP4cs8aKKMQWlt1Awt+a34c059ayF0P/tGnVEz4RzW5YuqwA0stPh0RjZ
eymFc08m9+qmBp3LlDBX8sRG9Q5J0SUO5eSWq5INmZFy68iNV3qfASnllH2kmhn2c+RISQyCgwTQ
DLSKPTIA8mYf1LXNvgMSAgY8XPQzVZi605rtW3jrKC0Ii1EDJBMWb/dg3a2ZCnYhsP6wXzCwnS5m
iWh8NlR1MIg7WiDMQMLw6cKqzCzSFIcr7Vf4O8zrYzdHMVtFkdj0sd0HMDC1uZoGcA0LBhSyC4z8
QEYuE77Zn3nwg7Hgd2k0aT05f1z33qTNdNlxjA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 102992)
`protect data_block
QF7ykNjdxj5wFiEJghXHznxEuQZgfa/v30NhiflZ48yjBSbAAcaLDySqQQx+thVmMUvZ1wG2e6xx
L2vhbd3tKJ5mlzW53NMbHmBu3el06pLenPfnEFTJmIlFiXKd8XHFIdvYfWOlH8ZgjPbExYx5PXPo
LlNhkI1vRwLmSxEhrVzYGqSs8ZgHw3s3I9H/RfTkJ81g6EPJEBS0eFNpyXtAAA/hTZlT37ntfTFq
sBxBd+nUyltrAlgu/Im9enl2LMYKrxPOWnuf8F0/luXX/jWCtp8KRSyuiQmvd4AyKq2lxyoE6mKE
o6AQ11lPGyqfALAP8slaOs6Km7xbSdRcEhVdcqPaUMIR6BwrtnpBZyPUg9f8Jb3/JrM1kj7Y/rQ5
H2orceWJ9KG5dwrJK/Rlokd5CAgQlpXfxh2fbPrf5W14fiL4ItBc2fRBtCxfqNmgY46xjV1y6SGH
i8YD+YxCtI/XUoZy5Ivqbgph75GkLfgaWwW/UarcLlxKipUBXhwxb8JZD5wKivw75REb/y4nMSLQ
pWUVbf0MRDq2jB78bYq/yZsQkAJ8UP8Opx1YjKrzd+z+sTt0co2Xyhj03djT2FeJ6c2QMBOobqMv
Zm+Hj9QalA2I6odzUix2cPnqYxsWamEcmF0kZdJ3tadhYAouhj819ZyngHkrhGioLqSBbPBLJwEY
bypPiY1+oDxz7gRfxFVpZwuq6hHDDHavvZ8Ps5mFQ+8jjh6+eHY4qrd7MVwgDVLMJfkYyH3gFuP7
vfuKEUHDvMrNOHr8OjjTtAgNepFgWG9xmO3kk0JF3SKd+nhs3PZ1xMZpgwbGaam7J7K28pD+ng2j
oMwdEMDOVcnTd/ngj09vg3wacaSYOW+wT5mxWI042mBMMAZXAmE3ukI79TQwl2J1kIomWMSFyXiG
jRUSH+u7X4sZ9J2GTgguTFuL1Tlb6aRKGB3w+58ZeuTtPfAY0V1BQwradWZ7xmrLh9kxXRe8PpQj
0N5GFN3D4ZpWeMzrZLClraImpX6Eha74+8wXmxLchu4LVm7Af7qAw7S6WuhyPexExs3uji0X2HKN
jR9/J9/d/uWBv8WBYVWETk0y1L7vlWw9feBwQdyaPlxkm5mC7oVGtlDzwGzJaUtHjFTe4pxJ/4Vx
o9n8b+RxlibghASRUsa7Bw57JwmZDkUf1ZYegGhvY31qZSyd1+gLixfvsf6PgWWvr8xAea3NlU7A
+un87WZy4FtWsSVtTkIObgw+UR62Vr9DSr1k/zUrsI7dN8AeN5Aw/fTk1zJIuhfbW47duW+WS1FK
GDwU/pFvgr7diLcmpxEXMqiyCk/WEw1EspTW9wFcvIT9Z63HSjunXwkaj/73Xmwq6qu5B95Uh+g9
o/g7TVH+gnHov4d3vbCPPbqJBiqykHB6GSd9U/3sEb7IOIW+6xFBOWQDHGM5KZLNIiXnbZPN3yZc
wsrv5TDRoGdS2KpIyjIvXtJ67WH6Z+CfHAxbNav8y20+Mig1CoDAqSUEMhMx09kYbS6Vqqikn5od
ZSot3gWfx1Y2Y1ncWApZdnO8BcjMzM7yMgm0TlX+EiAsLjMQyOCfF9xzskrd0OILDASVDyaWoe5S
XUmdnU95PSIJp9A8RXMmGSUCwJ4uGZ8xHi8tG+bf4zmYFNt8R5JbwoqIpaekLXIMmN8sgicHJhja
dNWjQPbi/D+DHdjLMvYv6ssxaz46joHe8hi/gzpwyKFHY9I36xlUcvBrR0meFNIBGn4EMhLIHXGC
yar43aYG4VMC+Fr5o4ZhgplLVqZyMTn3k/JlF78CXFJLVnhXB/Lo46Hl5eyE3ioZxdzKsg8u2W7I
D6+d7QSQ7bjKFKBxBRtUv37BqzhQwmy39wUjOIukkjMbFpW4PZjjyArH4bOxx978Xgz8ITgMxbFs
6KdCkwcrVzNvNXjfLfGm8W+IFMtKX1Xxrs/HkIdcGIwCrSyTyZIeGvglv0EiRHuJFUTfUu+8fBRV
nOxAhVMLuXrW3MwmqV5tu9WnB4hJ6UYcwpPVbeJ08vk3bYFUNp/wStHkmHHeG+oTf84NMCSjw9to
u9HH6pTH9lx8h8zgfkuSblBKdwNt3RWDF2qYgbghhL6dvq33hdlGo/S+D7xjgz13E4V5EcE1bkxP
d2OHtRT2mxsAWG/1aPD3soXjJ027/YLtEfK4vPNB2U9kG6F3ATPclkRb/WFxfDIO34NJ9oypKpJs
tS9SWZTfgVldk9bt18T45ePvFzN1Oxfwv0ZKOu1aBqU4ssBoO+Geub+2imGhVxHMVsAlGhfJs0wu
DObfDjDW0d35IV5zAdn1GH9PGPHAQqVvmki/azh5pwILbSejYeixrBSl9UllwPFymgJ0bFZexshA
uzY+9u9rsDkm+wzDCrd2nvw2Nj+W2c2lbkqYKwYlTqawrPDHN61pr+M4+29siSPD/3rzs2dSJ4m8
64hIzQVPJLIKOfT2bPuA+sOoLmjUeOAvctZC5YZWz6DUJ6iFnkoMIfxVFbyKfAQhij3ECcm/ccSn
3rRZk7H7WY9PBtGQu77fVr/21Jvb2kY9feugTpHfkXvrx8e6zAJJgMOlRhs+TNhAkaU+mNmLTuRw
OIKAGQs+2SZ76lz1mW3aCP8i6/e6L1oQgzDzWsh7WiYSKoN9ez9Giekw8ZWIXSCVM32P9lKUFuRt
ji5Zuz2NnqsN1Vfvca4pxhcTc2T29SoI4mwf237nwHaTz+q6PHP/Zsyrbod2jFDLnymYWRp2lPZA
+ig77kcie4v40JtBzevlIRUgMM5YmrW8jIfTUvJiiKYj81h1fhU94Vh95F1ovYXyvkaKroB1GLoH
TDYjP+SYooUGgqK1ENxLtK5WJH5zveMtWz31X0GQvjjz/hoBkfmfrzORyifrOg7+Cdq210CGe0hE
7Uw5xbyf6wgjGVJ7DqeDaKrqDxQCu9lJA+oRYQNDffHbr01Y46s8zb1AX1b1Me3cMwtZAtaPqN/q
23YX2VgFR8qyRYawB6TQZYJH22mxD1t/15DirYbuUeE+gRHYPsTn0nxOF1lcJ2OYcyFFM9q87EZg
FV8w4wcK+Az4OV7F4Dk2n9puKDWxAEoZ/xpGWwhR5cw9dJjayDIsctxB0f+8LFgmMBcufnRlXgs9
Nd1EWDYRSgpFAPjmY42N/Vt2QezH4TBe4OXAY5Zb+9Q1hjobdKlsHpHLCExN8sWce8peXFfTDPpg
9WPyPOqQ0vhQUJ6R/G439YIRIG88/Yf0EU7Iga9jTwZqf9YyRdnzZwqoR5MAHLBzF8FdecSRmWkP
5tEGVxgj7Jcsl3csEr4KEJr/FgAtD6Y2KcUwu2gXswc1/7cIScfyytDf4pkBGvsIM4I4onfQDmXl
Iq0Yqlp1dtRw2eEQyc4zhwzmi6OqE2QnvDprfaXg895F0XIA7+rwJr3o98KIIXzySWJNn+wnlidS
kMTwk9sulXIpoqrMGE17xQPeiHky9n/9MK/5EhWQ8nfc75zn9Vjrw1COuZRvvxLJY+CBs8AU0NoH
wPTO5C8bRThSomfdti3Xh2ASLXwy2606zn+0NkmCR6Qk8dxN1ij7VhAyz8UzRJI3QKAKZHMBdzcp
n+cfIXExn37CfQZYyBp2+hSE4lJ49+ssklQQ55Y/WM35VDIRCclJkfQKJEGipM20ulD2pUMSBIB0
xlHTYHWAfMPiLccJ5yFYaRSHWmjqE2K0ODfqCRm9c6I7r+ZWH4fWLyWqsdmWfv3Vmfqt4bePfCfV
1fXerigdKhm+47yMzoB2EzTvo+cmzJN9ofJlyv4lgw0f9aDTJbFs/mi7tM4/aAL80FQBjX+BGNXE
QKi8aEVqPFr4MuwQMcB6Ecisn59GZ1a990AGC4tkZP2KsNHLMvGxDqv7WCbDXTFuCbNar7zVDgvR
MamzHayvmnss8ZFQ4xaWN3eyMpyE54c791RW8ww1Ld0jZC7/9umy2Fa0mtH+kBTjpQu3zXjLAAji
6gdzGU26sE4Fht8kWjc1Wn114kTnlw6CUVYZYF09CtBaghEL6dSKri8KgFMWR/J+f6tmx5X6lmui
Ecjya9JFOzBG73SlLEq4/5T9BIpNSxWBJfdVuVB1n4QD0h2cHxcILV6wsCGQ6vyXc9SdEAtSp7Nf
iXPqIrIHjTLZv3hMU/MtzrBs0hY0FFwcIyTRgQoKhvxVgHGUOdTsyJrELCzSaUs+ZhOwPeWEzuN9
Ywt3bMu2FyX/CNFarDM4N2Vz0+aaZUVr9IwplXfJYrJJGSpFr//X7CssVSqkn2CSbejKHe4e5YC6
q6M4ZOsX8bit0O3/EF0F+3MHfv2/AwFP3SAD+UXYD0S3RlV9nq7rcYxFEiibJRu6zzN7SuX1m8jl
qONw6KZobXpdh1l3Kv66JcE3Iawef0+hhDz4WLd1iI45sRxBqFa49xblDlrgQjmZ7N4Qw0v/SPgL
Y06qYgp9UAIKjLw9UG6XjvGbWgm3XKRbdzhe0vX7DQul01g9YGX5AIPFQc+5jdAMHBrLzerO35Z/
BVzD6E/K+ywtzNKWTnkF0mMoBsJBUAhro8tj9rWs/WndQIEYVjOKJzV0dHYXk1WjGl02eSQHlhKK
fuB9MErvpMhRfUcB5msvCNl2YoPklktt6iToT0EMLzbZiW9uPQ0ZX48YYYwF3IUQZ0EwaVdE+rqo
5ST90HR2tHAkjMmMm7PUDK0rt54hr8jHqt7+VQ+GUaomkt6kaTA/5dgpsksz/M54vvAfNdyD4kMZ
ixoLDMpGWpLO9h4m25wslIqeYdfOmQlKM3AfrSo0uV7ztW+xOF+VckiyO+3ZNhHNsovMH0ZajQH8
ijVWePP72VanzKvIVHSA/c4fpxUJdhDsQPehVY3pKgwvsVLkROYo3GMUVMUjHCJBEq1lqEbFRSTG
EjoX0hIO3JsL3j09dLNHwoTGrR4SUHfCllDka74Ypuz8wILymaF6XdCEzf0kayoN4UISepk8PwFG
xsAlWUNJEvxthhWXeuJ3GCHeYNETiJYDw4jHWn5fUDXzrQdoH6v+HEUiHiP764GNfUdStcQF22bM
KllSPsvHHxFfRS6TdQlfTQ67m4KZGbSLe0RXgkGxlTlYKT43n9rBaLDzvXmbV4O06GC1CMBWCN+d
g9BPfpEI0rtKk0bMRP7hnx3boP1ChU+hsCFyhUK1VYXf0lJV2fCXzJda0hVQBsPC2eFyvfCUugIO
VBl+UN1RmvW1n/+ENM1XE0m4SvhYIvoLq7RrBYTJmAwNwO52pP74A1uROQPSa5EmBdlKnQD9h9mU
8Eis5piC3QL4X7lWRtxzZSJTfGpBX/db2H3Qi7/ZxAppQp6s1x2H3YBB2KCVd8hX5lmtQ3gBaGj/
9U/N3mjg//18Zsln7SYmtDGxt/wZheKIW5L8hhge9pNGw1GE1qfZOXDFVCBCjDN6BMJIkQSql7G7
va4AvSt2SdEIACv/LioYf9JK8Z4vm8l6gU/gVF3evaaH33TISE4KgZ/KcKQVssMBUlut/peOpkDr
T6dcU40R/gl32mBRlNkpoV4zvxsvh9KGEBuCo5koa0ZyFOQdC+CT/4L7Guiaisj1VFN2cbJaaSQ0
Qsfa96fNNTYWG1PMKZt5PXU9DrWNRvspibbDuYIwfK1loxajONi2k5oOkwoETTPjurChfFqeu1ut
mUJuq+GccQ7juGXBiw9M38O/r6BKFLp5fIRI0po1TqqeFL2AWmuVnkOyf/VhrZqWdCmbeSOb9MA0
aM8XsKzsG6ZFCsCUrSUWe+4JC/PjXtV4QSb7bduC535RUyE7Gh6Ioix1QTw4uv5Wtlzp0sAZ2QvA
8FWbWTJIQcmbd9xMTXUhot0RSpFCeT+4luk4I62WnvrwY6Hk0Y58WOm4oTyZ6U8cwlQh0Ty7Fib+
0nbdGPWldwGiCdTyNEcLX1ZyWizIGJCabDrzKu3poO3No/4Y86Z6Az6pKoDO0sto/ObEWISIFpGe
IjtbhrQmN/57PL5MYYDbQKx0gqYlSYZDh58tkJF7yPnPQJr/Tgqx7Uz98SJNtVB+FFOm19P+/XIp
gVLXZ9uKbE6EqPiImM8wpUL3ertaqm6ewyAEa8U9ezaoT+CEkyogX5RVgHRXOhuNgfFU85vyQZ2+
b482KvHoDa2EHR45iHiM33Aja7e/mdylNflnRXNdravkBQpC2jkjErBcblphLz3P6KuStwRcTnxQ
L6IN8RJQWOi3ZuXUGG32+C3si3cyTN7tdtL/7HSJODqHOF2FR20I8tRzqcTBUKHrHVTzf4CFiBg7
CvZ2V7/hJP7ePQS0cWAA56U45lLzLSvj/tB4YC/9FQ1v7gHEZLW6Y4YEKx3S2ORR+sgzfcUaVHTS
j6VukHmEzNP378fw2dfjFOmk7pj5sKus/OHZcEjxqpdkph1owbNJZjA9DajA1TbcnagG9HiR+ZTU
bUPv6EPL1xcJmnZ/aulVGfXYTeArstrzzCDij8WEQiCany3F09Ph2hR1XPr+RKRrMnEtSceGPhpw
SyNKc9LZ6YsTexCgrLCx0TSF9cPyKhzGdsrCxWpOC0h4JPA6aOjMXL1b7jXu9vcS13DPqsdI1pfY
qvly6UFziNPShehtlXGa+S3y5Jxvq5Y3mYCgvao2yMoygLr6g4+Mu9CZ8wOn9yofvtr82X+1N6Nh
Fn5MoPlmKBPgdnXGBqIq5Z1WAM+9OddNLVFUMbApJBG/vwke/X2oQwhITJ4IpeEe7GmC9K08iWZ7
soj8CHTEUcco+uUZyAM8Hp7r6hm+3FHsZof0wI8KX0go4k0ce5M2QU5+8uQaGdyQ78pZ2/bMTm6N
NmcRZ//UtPbfSjYqX5JvdlstAw/NW4f++lSBThDC8y8TCKRAd5VCGQYPK2wsEGYczb/WbXcwM9Tk
H3lPIw97CVH1YFKtwnHU+r5vVPn7fwS0eEzD9xqN3xMLsYJyylkNVwRmY1jips8yt42K7zfeJHTX
JxzKcNdBUusRsYsUrLDwZpoFYRK6RkEAuJ7EQQun6YQoV/n4CeefPjHnEcKwBFL9w6bVI2gBfmQk
DPuyj2kbale1smyb/PUjK0T62FadUnkqgFOkrBD98GjDnbWE57QRZ/3keFUCrC1/VWEhtn/yDRx2
dxI57NK7wpiLc6gBNeuU2uEyDetzyDdYCfZrdBwqWx5Ab3bJK+mdqEhQPTVbuk1F+RYHKivnMCHt
mMtmfTuF4PGMV7t7CpaXG6AzlmdSq7hCS42qYxVO/vMSFenZtVNr1JTNhDvvdSsqIKi4NZgi4+KT
fMQXgWU1pSIIkKuoAStho6cVh1N72v/fVUFSMzXdmYMm3msJKbXGQXb6F6B+LF7HVKMXcl3qgGid
0b3m1QBWVr8n7G/1mId7CLPsztxp3PgqV5wZ3fpiOLJe3EbeQ49wY+2MONs2zO/+GzRENMF1pv17
4zsm/02veWmTEmC3v6zg/eXkTDvUjxoByyB4JJ0p9bqYgUUeV6ZH5hBunK/bJA8Adn95ltlSqfrR
j/i876Cpgcv8Ei0rG/keDtmDD3tIqvolulKe3s+nKRJQbQxWGtfuc+SrP62iE6bjlw6mrFaadqAS
adaiRsBxhMAJuhVlzJBMrw7X0h/+jgmIE9HCZJ2ReMs6uCrn66PkhSThaI7pR5j/c6VadjOiDfhu
FcGY9yLXaertMnkBclPX5KCjd8+lRF9lpzhFXQ92vywxizf1CjFBYLLTnPU4rYLgy5tvAkm1NAD+
okvi4Q6PzRmPyuhIFFED84mgj6eIabvEPj/EaJsQWifKm3sfuPsVbz42pigiTyNejYrIaekLXvDS
NfojqQJtJeqnotiKAl74AxjAAC7ny4z3Jsx586WYDRfxG1+F+UsJoRfb2IjLZ92p/pIG4beMPLx2
8YnUx2CWZFdX3W+0F9vkMMx2x83NSIxkaNeBAHqFsH7RQ/sqDLluHPMfrjQqDkcIGhH1zmOlc+tM
MHQb2Fkq4BrYShKEycY3F9VE6KJj+XiFLANcQMSeL/1RVAMwS0gXaWfmenV1f3QNOXY9YuULOdnS
96o6MMSIGhrFA+wjIk+GBTAc+prLoRhRX51tNr8Js3o14BxUH0ning+WQqA8Tk5PooEgXbcMpumy
rr+GdvQv35ZMc1O4xJ1T9SdBJWjDkXrlfoOpsnSIXvIawgqcUepO+QKd4QWj9MRrWc6fFFrdei7K
os5S9vX05Hk3aBmASqyQnnPC50BqJQwx4QqaWmA+yZbJq33T467/lRS7AYOIpe7/YKSwAIwI3xq5
qRne3siswLVuv75go18wgJVAtOGfSUHO/zFtjx8EIehmM4oSER8c/vCClpg0AFPcmZrPwVtg8agX
HOGDJeRjffPfsRhFvvVmVQoeLY8J+3dfFVT2cow0DGbgcmMTC27N22KALShXiwFAY5aijmBXZmQq
mOjSlY8/ap7qzgdM6H1uixPXzaJ+dTqfQSTvbGZudwzsktpsLyuMj3clrnHfc8L9/GIplB4jiu4j
7Gt8/vMkdgy36TBqnhd+8FDEYZmfgrL36PUbqDG4s/28Ss1wwLrHP40Pkqm6bLtmt2JiDvEkrldz
gmm6bM/RrUjzRS8hnlU5ZRusYhsg3oyXKGtb12V42+e0UAG5v8tKfdI1JxRsnYAg8sgLjLGXeu/V
BZH1t5V+DoLW5h/HyQxaF+kpzcvSCAHW2Rsw8mpfVAY8u2BUW24XM9IdX7xoGHRON9D+X5t9z4fD
j+vMywlPGZH/HoMNISRYR5/K1Tdigp22iJJmyIsojQfeZ9+a540ZimhB8gMtYbkzoiqhrP7+Q+hY
8xnO8v43kVG0EAZMHQsfjP4tJyKKEWikaS9V0JRicDamrW97PqnHYMSBmbYVCOJ0LLHn+NnSNwdQ
fQcQDAhn9sQ998qWDRM9Hn2vxKGGxxB18sbIPukpStM9UJtORdxTzbqpHqOBMiZ6MF0El9zbJ9Yb
6iyiVe0NRzsGGezqf6FDa2gF5TehgG/eHQs1zSXvYzezmtt+rOSPARplmUzJrHrQU/iaqyQE/NSl
PdcjKvG3MqoogNwky1DVSKWDBc2PSoIOuICeOrWlI/UWwcMZ1cmDHg/N2eBY8xRZmSFqQd7UoXT6
UdrZz6qJogFVqqj8zEKHzA378/fGFQTQ0YQkVZrYNmbNdI2ovmuUByghwNGuLwiFe46tJix1TrUs
p/8MRIHOF367W/brfSn091DqIRkdZNSSkKGUWQChwUcrC+EZdpCdAEUDQDjLU+x3ZzADrMlMMRmS
84ZSQn5lm98KOVxzaX7mhCQ1DOZGW67xpVoY2epIXAtzB70kPVTBf8odjYqlxYFzZ54GIBb5t7TZ
ywcnajfbq2GXPVInjoo8NMSfxwdwyh5NpqPQ/yD9pxKtKITdkJRoN22Xq6taaaWVzi6/bSNByiUe
BpOj03AaKgxUXA3YVxKbPk1ayV8mqZUpq6zFu+uI/6J22lQzVTbZtHIQwVCTdyJZydnOulLGeWI3
Agf+N/Lkkh4fm7HYWXNMuXF5tbi9nUvBqUMn5pgo1I9uKxjW/pK3LrSJl7vY1HxG7nWpQiPa377U
DcUGuQ9X5VyaubcwQ2dvMVl6vSdVbIgHTd3x5h8Zwj3hHdBeq5HUBSWEjbLX9QwbtwsF3eUkN4zO
w3DDEGkeIiAElC+32G32pOT5ZZxGce1fktz+3n/9maXH7bF6I1A30WHG485sd4azcqQx88rx41h6
JJXO0dbDQYkSO2GMeeEElaujrSdyLrRASlj803z50O5ptdKFuZGCiwjf76u4c2WSmuci9kC3Z5Rg
8IjKk5J+7LNGQ6kyIGlNtr9200aWTKIbyXUyUL4aJZ42JShcK3nxaSflBraVYmO3Hvg1te/65iVp
WFG2o5idtfo1B4btWT7LutN7W2TydjI9tbYHEQmLBehhIQ+NdvfVnfPMiQbsMZ7dXBtHzje51bMA
hvHPXjaHjYcNEUNpZj1sm5L71t1fyvhukqqbX8vYkZj9QEJh6oLf1+a4YTfjbaMGPvIjIXE4krzg
NUrJE0/39ii9gWXT4oHm0qYugedoA+7KiCN6viiu/gNIpHMsmOLHWwRGRO5NpWgnAmg/5ykM8w9I
mVsYiVmRmaysqkRLNnXMkV88H3V2/jcmTjw7d0ijOj1OlSKv/LZzrxEiL/0pE9AEIZOOqCrSX4GQ
OIGURYN7PQ0mNS+tir/MEGa2s6yecP5q5kKyA3FWYUPmMR4L8k+r+NAaMZ4cCfnjF4ufHZ8UmvBJ
l/IzP3RLtNjuObxcpuNYR1Njkubwy/m4JdOtYlHbunEJcNmk6SQpRsWUUMq3UJH2gWKZ17rL8pDY
EA2+d7OfCTPxv1lib5FA1JxXwGGDcK6Hr42zQz12ySeny2jZnGj/I7nS3P+ra4b75JljOWKGBdzQ
nSVo6/tBpIBHXu6b8hY/Gi2/lr/aEGeQJPJf/Do9I637EJj+FiCk1SKGzQBylZbAEEbuJuKrEMew
fzaiCwBJV4oPzPkJaQRA0d0KkWw8KwCJRX5dIsKX0mCAsemrn0yMNM8HCYyJD3KSks0og/KBHBBm
cvWV8dXZ89MLw4JMu2sxR2xxJEK8KqSBeLXm+dJRNJ+ZEgyCfnVKS1zlE7L57W4nk0UM9IdR7UEm
BcWHZl/GoqjyM/plYONmj2eRFNgU/mYxn0A3/95RKx1DB/hsyKJNko6J9lPqEwNZN9yZ71z7OSRX
gQ440VndjKL3BNitlO89jsno5JSqaYMuQgXMLopU1qbSlBALWZOug/68RGi2JD2/+mWmmgvGhYuH
kz7QPCfzIZ7SK/IisVzOVcckSC3SE5QNDp/UV8+wnVELh0BSNtyQB2dhj3uPCkLFcsbdCkqPfApz
dEeNvZIxa1d69J9szpeDwe0G7z0NXPUTeOs7jR48tMa6Daqiwl2SOG+wuyPolL2JTywRtzCN5K/+
okAGTF5IvDbWCXcRniHZ3opxN/a/lgChfoVTMUkCqh6LhAwo2rtIbrGctS2z2fnHBUZd+xgF4beJ
K7MBwSz63C2FK9u6MwNT07jX1e1rebyb962f6WaRb51Sudy4eGITWGI7sLz/4nsqC6+hWT++gAsK
BjtDGA1kzkdrYWW78fjKrirn0UBwCfhbHvd7scndBDQsdcmdXr9EGVndPxJTDoSODy1PnMOmRZfR
PzvxnLqbuxKpPdCrQr4A8BGghiWxdVJrd3CCWFqz4wZojhoBHB4XTyE5oxGWCWW5lL7UX4SV7IED
n+czOFTLZzFEP6a7E41qbr2WAHLW8dA7ZHTr5RMxxVwApoiVjuz/TIia0NgAyckApgib79jS/84E
ctY2v0M6I44ihxsom0XaVz4pQZbUWXlH1FPLQfFEsCK+tX+Gr97fjtIZsKWOoWn5NDcs7nhXUXHi
3SUbqCnUCv7Nyav9OSwO978k6LiEDA93uyrqtAQBj5OKysj+LzMuMGmRpyb87ETbusCt7MTbYbHe
FmheTfo6nDEjw6E/jXydJ+UhT/ppplkDA59k0Ic8KWW19jKT54wZDYFyCQRLBb4+yX1zN/hJqAjp
FH3+GCEUIGyhe3H9RR5gjxNJoNRaEf5cFXOtINc95ZaMkNn0jlzm9Ny6ndU/oHkBlwMLUFtZV4G4
9+SRsAsWV3E6D8EQiZrsgYOqVm/a7lDR3VcrS31iksYXowhFV1fBAnVVC7NydsrfwyHtw5MItxSZ
s1cXFIfv/sl6uKGg/JvhSiTFR4W28nUC7LhVjI0s1wQG5/iQh5AOojudMx4v21LvEkGFrkY1t0pA
dLa/rzmAgJiS75Aa7QUzjyO6xOIaRisjf7pFx0F4YvR87Ynbq1Jdj0J/U4o073moxNiwEzMJWmNH
b40bwxuLK3R7+864DHbBaJjDMxqbZhx7h9QJR5rMfFoAk0LfE3AmcrLeHjnkGTdbleNa3Imvoin0
UPdSKr7jWsEe363N0kN2JsIWm6mue2/fq/5TaKd2Q772bxImhgWIxcnyBNkaWYVp2iufHoCo52Sh
Aa1VA0DeZTD6qr+ftqWfgFx87Hdmdri0bvCjT7aAO+FNkxe21X6STay2y4HIHeEDIBSDfBRfsdcV
ZGUSkoCGaLkXIkuvl98ljZf5X80U+5JDGVCoE39jhiv/z1UOJnWeiI28avFcKUaHMY8Xs4NnMU1g
u5TMKDYUSsJ7aFzcW0BhfzudgQVDOGMh6GyNkN8u5RtsOfrx1nnhUCGkM4qgZRl41g2oBL9/GHHx
lyVTOU2anffG1WNRyJ/0fJLFpUf5SCUFuGOplEYLIDofXl//o5FcGRD5nMFJ5tzT+uDh9mAa2rVU
XoaafgNJ4/R1xcVaLvjymc1mqNlmFcbCwwNzZyOXPvI4tnyyvCr9LvWwg4TMrBwKv0iW7TrxtGSA
JjlFrxKZiNZDxNUOoqySw+y6sEBdjLnm0rPYSZ9FBBw2lnV0+NgRgSrYAgbeBs6ssr66/4Xq1lOs
BkbF983zKmDa1EGBsZPFSQGxZ2udVQMVKn9lXplksJHBfJhYwDirIgmepVhxeX6kzeIlcHBGvX3e
lR8ST9NuIgm9oh1Zkpc6FIK0AJ49oWcug5S11B1PLAXae/a6gGXiX1S9Vc+0xH6F8VicCp5N1jIt
xz0PSsNyqnE4Y/KvzeinlMWwYXc2gOYCcFojlvIKfU8J2wuaS8BUcULyCQZRhSQyhlPx2pQVBrHC
OjgYcN5ESc2RqUR9ViOi2K01hNi22ojj5963cwcxzdwv0PQcOEr4Z7QMp3iZ6j9OzW3m5pA5jdZG
t009CjtIGgI0bulc81kBsSv8qeJKBNeSjC0h1+4PK6gWWarrM+DgeQZ3vkWcgc7U18U8G7795Z+e
bsyXEPrfF9P6MCSZSng18udxgllTWXvsjLxLVXAUfLTBmUriggdrgNWqCvEJwA5x3vVzLenZhrqr
ZIUScsfykCAl5xQcdKLEsG/dCwfPoQU/Vvi02uPtsQXxwHoZGYa+dR2kRNIMJzaPC0en2sm9BZSJ
TiG6F4DcErWrWWQSreemKHlZtcDQkqQ4QQOFONXUPkh8rz8mcKZ5bNS780iiKKieeE9I4su9knJA
nFP1ov+wQA4AQramHXrQJ2SBI0RutcomFkjv4dXBuEIoYmYIIQTqiUoommJ6nT/DffAwqnMcoISw
O8AjXQalUj+pWu2U7/tEUhudZB+hEn39mN4kIczoRtqzubGxZZfrXHqixhD3GCFOu+gocOP50jgi
PhAzNcOV8an2pFTL8s6LtaqYFT6qaXcdywGFgp5Ih31hfhwaTDXixLEdkGKBJ3SYFzd8qatwD1Hx
tT1HYP8GCGxO0iiwFhc7OSubddqCrc6Qclu6tlxkORX8suVv8YP65vKSflpKF5BKdzd+0CPfBEp5
Swa6uSxGgeM1Arqa1flcCWPDNWg1HBuM/RznXhM1sDq2Ve73wOJlEArwz9HwxOTGjG9mWZWlwXtY
tXm41OvQbxT3Jg45ccTAgy10RGGFSjc3wPZhg9Ljt+ROjMxR/LW1ZZaT6lCv6D6sta0QEC63+Tqw
tcMraYD9S4S7UWld+6eVst5z1QW0nUgO8dIzNeqetkngYkNqaQPDo9tftDXMoOR0Z2icUkx1oqFA
ZTvKgm9vOfoA4NZj4EPjfBvrYDBuRr+RHoUChof2tDHzc5S7N/wHfodhO315Q6TE1/kGyHBscp6K
q/zE2EEM6zilBCjdkevl6bxPvWSUEEqPaQYrZi2DR2qro9Q11CqeGzum3O8IIohqDdHrAIbQ/rI7
3w8SVGnTzI1DctdCC1/UwkOg/YSGFJd7xoe4jq98oe37A04lLbkWPVJX04FoDzUm05zgAciD1k2u
Oe9ASahUSNYvGzVoeJzB4cFW/QYmMOjKccdX0TR0B9lWPPhDKiTpfPHeX9S0pMa4HVD0sGrkUMPg
gn5v+6zE4eO75q5fQuW5eddCQYPcjmymrRQnx//hU8Tad/eefIXcY46hUnn/zpAClKvwhBGgYA2K
7XiknYIg8rum47kJ8UZoCvAoVcav0zJmW3wfGZ8GWIZbQRqT3gPcxMNYtPnZ9q7/l7b4t6a0Agp8
le+QdCyaAVk2U60wCDpZMpejMNOLkGGCOA2+5AO82Qrcb2mWVsOv6ylUMz7Va7f2bN5c0a2uKN0g
N17a/0jv7NJhFO63+XTxfN/ulIPUd/WV3kFEQoiBdAQHmxJPZ6/MdrLUbu/lUmZ2FxXoIoxQcuRs
2s5XFLNesJZCUYo5OspfZtHo8Lks869f6DmpyM9gIuFBGb9TUA/ZeheueI/jxQputYSdfZhJLeoO
UaaMrYITgpouXWjrwjVttf2W/pGYir0taN2S/nAPN3ILVzyjjJbDEChtTWn/LyXHq7R9mwgMiN7N
7ZCkEaIe1uMVtCUxmGB7VKBoispsiGuvuaXqoXn2FnuXHsJNQnv3zMO69suQK/veWnkLj/q+NX/H
CgjeBSlsPIPt9mM82cv3JJiBs7g3vU7yJDsB9V0nyJmsTYMEeJYTrdMvqI1feaEOZ+xNXn7crMcC
dhtPFYCYNY3L6iaX2Gc4LeQb3h4vFnSnEvhkVAyRzXpuuGSqkRMkGu3S0D3bOagYyshlY8vdlcOQ
H1RFV2fcCA4Z2kE0C4SfXEOu8DACeJRcy43EypB1iqRGakjl22g/2DJhssPUIYRuo8Pv5xdKBJvq
WKjtWBlBO99OAqSnyBuX767DQZ4BS4LTur3qOU/Sm1RovRaFn2QCjp9PPloTvKIH0vnamPqnvlmS
nLOHHNDegMs5Xcwj32F1m3ja1IHdDKyVLGmN4xZ6rMWvkcV8cXYbVoFxKSqrONK8e291+Xb73Prw
94hQNwXzn3FjzK6QnwvZfTWajhfGJeGtYLpy/wK6koF/QyWMXfbEfXdt+Y3V3IUxi3nW1bCCcx67
8wsqlaeoooDa4WftxglsPRisisQJCiGVuIdsnRJI7Bn0kzXZBPkUnUjro65nEpk9xLEtFYgAbyJ2
tO9NxVsZ8LGqFORf25ZRmrWK8cavTY+VTMf8Ee7RIOBqzI24ETs70hYJ0fVHhHBPfI/tEbvDQm8v
KQTIQBjukCYZTAuqzUj20igzZR0d25IN2SLbB5Prstk2/0EaQZxNY4Kk8DoHxFT7WNQh5QxBSCiF
KJviHsyQg0CuO3MmmbUAWCXAZMObKuP9JDJhQn9Dxjyjk9zqXfAZC39CqbScjEw13FbZQZ5lRqgs
TENo1CjXJOiRwwUhThD2agsLvaslt6obMH7+MQ9jthSP0sbLS8JI6kivRwSIZsuRoC7t/LSm5tX7
ix367oVzUFfanTGiDmf4uyakh3oD/sEd9uC4y6ESoN7XTgE9m4MSoRkLKzGptzge6wKg8guyRfk4
C4QHRmltL6FQRriDcRkMIv3nnQHM/Tq+Y/0aEbzq8uz1sL3uvS/SGLjkRRG2dWvK8Sf+byZEwjJ0
CPjjiVN9mOZeFdiDNHy0xFS4Mbs8K5PO/5ZVCPmXa/Tp/qmOfcMRN+0IwkikcBi//OdniJeeureh
BXMJsG1gOf8qkXyZZXu6UY+Lf/kZSWq4nrgWXL6uX2wUgYmyQtnxaPpOz0WuUDG2ZU3rT/A/WU6+
66yixlCzf7Qfy7/kXRk2fZcl6IQCYACiXWRg5In6wCCkTUnslzvUIkGHi7Q0O0HXCGfUkXlOCEvj
Q0VUudLqPg2r+DIZflyf8WeDlr/0H6sFmbbW8BYAnay+FoQnTNff6+2iGFepI4XwJu8hz0O2foN4
dg3L5Vektz2Ssx7XLuFrbOB0R/zr1Sx23N8UFYjToJLT8vBtV4ElTzAH31vKiawMrf0XceUaF4/Y
GLzPZwHtE43CKCET/qW+a/3dtnlzCyvYWdgIHd0Q10b4wpi9SPFUvuhmCcCpv5cTcMHM8AG5tXYV
YnvCXg/wmB0PBEhq9zOfHG2v61NJXi6oqNkHN3q0bYkwNQLjpT6w+PZnorRztlSnoTBGZRqbuUB+
9aYOi49T+wdD+vSCOy4qfEGUClDkA3xE5iv0rUhnenev7BY19ka3BoRF4G8apphPWZM91frY108Z
3h/wG0KQXFBrdkqB4br06+M2vHmYujRt1gQ6pYQuPT5JRLh87q9uqxPWsKG62ab3/iO7h9XZGKio
kRQO6BPdo6er6+jZt+NPe97A0Bc3a7Nkc8c+xUy7wnf70I9QaAWas8RuNA5aZqHOr6Yn5SU/qq9U
jWTKwcVg8l9BIz7k7ga03P/sucUJ3HZNMxMKC4gvfRhDcRoeCi0OCFgW2kK2Cpaf+VE2/GDC//gb
TIQD0kU86NsKfkV/a4BIkatYXiGNk6QNBWWdPd0kwoZ8vdie7sIPygjeIAxl9YDEF/PsTJO0VBbG
XsgAZ905wRlwH214vjHfKKL0cxFefLyfnc0C5MXWaL6NeUG38xxRmkJTvOGkCpP5ZO5ZQ/wIBCHF
6XCgLmHov49aIFkIthJeX2cdQj7XGdqMqbA7uXZXHO4cdhAjj/P43fr+zbU/1NTA/LstpAPsghBV
ozND2nKSwmFMvWUwNXsjOZLD6HByuHFb1DaSjnRt4fJ4F0q2K6YeSb3VJD0GwxZWUVNhFyPPGcdG
V2hdiq/P6F98A/iJTpnen0p0HugllYgov/JUxDKXE/B1ogI7D9My7CNUsiQDw6Wf/l+d9w8/Hcn1
xyPTfPnbuag3K2lGC/6uCmEa/WDEazIKmp43hY81A3TbW1HDYHnEHDxFSKgeg0WPg/Cpj6JLc3n0
7bfT115jGF1pBhjHf904skj0mBygP1mFFR6lhHoJrXXJPshswfO0AwCByEfqvC/305043I81FB+m
LbmriOOC9lhbuyb1l7cfIZ+UTxKhspF7JYh9UNFTI4TV2NyPNdaqtF4Y5LHfWsQzTr7DTnEkBpjG
4ohkeno/PFbeWdcohJehnQCtAiRq7NvPfCDG0VVZTCW1tBbsDtO8do5nGW1iRkzSivmuHkzvz3l4
d8um0TmXiB5OtHAbWH2mdyzBAsm281edZQXIVQb5jcWhArxfuG5IJZPnClsKb9yGx7x75lwCtxY1
i4e8c6+tTdQLI041ieVjL3Vj3q8+SGWzs4yw2YyABie2O7ii1Unsw5QgJ13tcBXzi+K0v64CgV9X
i2RqP8uCVX/FiS9jQ3nIlWZqsPcrNn37dlah0eqm5QEZXkG87lMtqfLysjnQDk8kkewh7vtlsnVw
M46vgeX5jnAOBKxJooHzccGEe4X/trfTrepcb9a/d2FWbh483TUIjp3SV0r6VjnIxcvez/NlHBte
XHKr3Obws704M5PQiqRn9nk2RqUbXb2FjoGEsmgPvizC4cyDd8sfEqH29AW4fKmd1dmcPaPRsm7j
T9Jot7g3FZZTzcKRbtxj0RMoo37bGxdh8fHf7z+zlJpwGUc30WdjpE3wR63oQeK3IB1tjRV89DCy
DywdWiRzkIJ47TSLsW5BnM7I8Ffl96kR/f1U07tbI8nwj9w6Uu2O6jlbi+O8ZiYTVorWM0G1NWrs
9G6/Qi52R251mbPQ6xcIAotkayz/HrsNtUCj3FQZoD1ndzIcDpMvAW0BeriWwZUNFhcn8F8DKc0s
oT09Gq4voDtz/OJRyzRf/4tg/O2iFgtB+M4XWeUtMSgDVIye78jiFatjvd8iJN3zeUItin7Uuya0
wRZxPB3r4/Ti/DnWUbOVXf7z9pjIZRyZ6XhkB62WCP7DsIO9K1rubIw1JEkS3hL7K3pfmkTFIclI
CVVL9NEEbhcmA03uPPIzIN6EBln+LjTl7qhWnlFmNYwg9QYKKlPNvpbrgzqIqfsdj1uXvxJHG9bC
yHQZOo2WxmsRAoB+YrvSdNtAqoGIel4nTPaIql8y0ilLnPf6SBYM3L5NfGF2wWpXtMF4cIZ6S0Pm
cfLIUtMyV0sB9HJLbJrCBKoBzSmCUwToNknpf8t4mW8iNqfaQmcd0KAd4tP+2WSs5TaG1ifkyC9C
j0Noa/2/i1OrKt+sTvZIa81kc1mKDGy5fsaRtHCy1r+XFWULuqjwD40Tqr1K8hm3QV3SB+ew+aEm
sRzXxUA0cjWy/Y8+upLhIOma85BC7s7M9swphsCJsrEwTp7qxNAaq4AmlFXxs3gu7IqfhyufTy4k
YzvZViez4Emi26TU/JQ+U63Ey1nmnOeAO7vu2NutB2W5k7XTWDyju3DVff/c1yvKXPV4PLnpvL5L
dSBKeqtzMKwEnXWKLzK2jlS1da2+wMbXZmw2yDW5EgECQ4yYY7fsf2YcgZJXN/WKE6tUKBWGuGnU
ihO4KvRY0kU3CsjESiVo+sU7OLio4xqUJJuxOVZA2t2X7e1vGyAQk4Nldj3qDvuU8iH6Rh3xPh5n
ye2o+U6pvH/A497nCbgv05ZmTRuEirB52oBHaL/UHjQPIf/BZg3sIlWvmEoUZCdYqxMhR5J/I4Hh
umPYxuvEreuo8VF9oKCARYPcD81EcFuIx2qkwqaRTaEcHs71uMh79E6Z9oioz9WAglprZ7AzsScU
/tZX0vDcjnuezb9Mf1tBZUn7HoKHzTRz/HLAKnumfMzx0C23uJ/cgO9qSn37RcgqlsiKjWzQiFHw
UAsiBNUowYquLFRVbkOsx3frRrPaEn/tuyVqYcaeeq6eScExQHqlwZZdjdtepHNlaq7yVHyn/aqH
lmaSTvGsSS43tyl7y0ZwznMH6ABgAR4DCRJC1oV3dFi8rnrQNwOCGyGWo1OTvHt5BMC7revPLPrS
jgmCaomxh4Dy8fUkE/mfNCXIofIyF/uIaGFE9ZqajtklWwJ0QNE1UPvEoIzLQct7cavirM1WRJMg
IVAG4ELnTr0tEAhY5a1a3VOxxxAosKwluL2JLwi+aOXdqFcr6Ya2/Q6bXMXSQucKnJ3kMkdiRaLy
Oc+Kth5SCDFhvr97vO9W/Xi8evz6du8lvetGyGe3YoSV0e96YPPqaZ2niAiYQnyPAgpaFFEWJ0oT
vMicUZ15FHhMVO+3z0zTmXU/+kf/4iTtH3WaQyjMjILuplO1/LvAWpHD/A+dkgOAva/EoZciKrOc
hlmvJ1M/AXah+8QS3ib/t7loSJxewUwRqoqcBD5bu7CKkIBYyexsy62ugPG6QHs/aD4XugrdHHsw
B8NOTK6vYDtDYVfO3/NJrEBAVw+brPUIS2dXo2Ivc+t+tOWnBfjb5s8GRxQyZI/oO0S1kR/iJb+G
NNdlCoqa1BKNQNnFwzXzT+lgRol3hNPPoeo+kqByNcPKR3J/I9u7/jJrYaC/SNyBYHH7GyihojBl
fi7Ob4PBCWZUhZFIh706Eg5KiVKmU0axrwQdBDMEmCIKSmhzpeMbA3syIti2wcql3/FcJ533qAEB
wum3XXujrYKzh0c7i474E+YHfb9BJw/kqd8e9Z0VGFRv94X/OUQXFjq22Ixa13rfokMNYjxR1Izk
BfDrk8JbTSwerzv3SUbBL+aeF1pIcaESRmKehT02nng2tWOfEfOrV3/Bxg9sIOaeOvpCJg+sZ7OM
KMZnvQUb52wKiO+y8bS8KUOPV8noBPkCwgpuUs/e5x6YDb9dKLVy6OpMfXv5WoS3243UZNQCxFF0
TG4O7rtQB745onCG/UxVQRsOAqsMTtYm1VALPMJG5kooqnqWV89mQlc6jiwHvxOITkQvUCM35XgT
eOcAlmbMYmD/spNrzJevTardrbk2IizBCI1tED5Zd2viJl1ZcpPljWiNnPnsyxdpPp8LfTJHfc8x
DwAa8JofwVFlIZlNtoQ5Iq+EiI45MII+YVq8wDke3azBs4H7m7E6n65n1/ZkQr9I/TBrt3WQMuuV
Fp+dc4ivv/Nw+p9lK24YwqakTxXz3KdBkg2eoDNIcy8tqMHuSsYvtiP+gTGx6VPMAZmH47amKu0C
ZMTdtXhutEVpeP2UjWAVHST19fOTlzZflRvXXwGd3ip5w9XhAtcJ25RL8XO9uFXdmYQr5YfcjIKJ
0dVu2K6Z7dcmZEXO/qf/g9sUNOY/hzbiyOOqdtzGqRdzlnoEpijJLCBCCsJsncCoNmk2qzupDfbh
IoHzn3BZP459yytUPbmRtit1RYt3ZTia7G/u+I9Wk5wf08t6PeI5L75mNfC44fL22uMXdOHXaZI1
Q/ke/CczbDxZQKq5Tjgmxv9lQtOEEXaVcZN+5GdHajOJP6tw++IGHCoJPZBxzpp/O3Dk9E7sNo6N
cv1xLQy6y2pWiaWjiteaqBQaJPqRr1ZItn6UYwmapxsLxm6M2pVV5SCYBpCc08wPu+Ok+UX3GZAx
kbMBRr6PjwUmesSbAJPlMHWMUYkRP7xIA0zqCha38gk/2es9dpqmuxE14CNr7Okm7fqFXV9UOCk/
EVsbdUAcOyLSRA0nGeyOPHo2nsh5EBFJZhr/cJLL+UPk8SEfoODpdjIHf6swrC3+O9NebNs7g9hp
E9RtWZvklicfnpIO2/fozjNc2Bq9jDz0BjyUe3+tblQICnVL+J98QBab6zZgtCp6YpsZuIJMSy27
hFjsrCOz71sY4R2a1VX8Q0IFzYHdRBkhI/yPSB91ycD0Y7lJxXSiYwgHd+xYzdDfDUnWh61QuqSF
M0vJ71JSglMudWrI9paE+UDwO/Hxe5wh3oitjHfq1+mTjyk5pp3AN1SnKD+rSsC6gWJpLtSOFfI9
li1T3qnGsNqITU4W0SwvzoB2OF7YiKni99fUTNJp+XaI2PPPYPSJX/2QbyKsoj/qnEGpl6od9/LE
twdd+H6YBRkYi0Vuyy4ATgtQzFpcSO5b4rj9TvPVdGle7EYZl1mW/ks/Nq8+mEH+vj30k3mjvaM0
BVmNqh+oQGHvlFeP6TxNFGQcbSD2K6WVNaJFKQ/TZiIOmFwr1eZdthEbiRyeuSah2Dwrqp9PlDyf
jJaLXahFJN+oM35zxKI3nZKD3P9cq+7/AhwDfZng8fCjlAp0jDzizXs1plvcwb55PBa2Pva38psa
razmkdNyKC9NDqZEMPIejtMsZ43PfC6h1QnwUu8Lu74NC3VdQ3rny/U5eA0J3YzweeZubK660On7
d1p97spw+pvkiBkgGvcmQInsBCk9vTqbqeKB6bTZ7BU/TIBRg7mVr0p4xWLXURXc3Quv4ohsFDNX
Mpmv3UVrV5Lw3rMrfSa6LI6SXIahm90uYspl/5FGva1hSLUijM7d30ECG/IF1k0axlyteNalpcUk
eT1KILC0//r98Lng8I1z+I1iib5oTvQgPTDlsOuyPkAq5ujNOL2z4n+GE8/k1d9JhKTY9r2JwgJY
hl3DcmihwZJe6BSkV9ysSSFJD+nmYDJeb0hCpEWlOCE1GnC1iFjKUId9y7ElsYUd3d27MfyA53fN
rIimU4tTFscwbyXaQgXGpEF9q5lIgfrauI+lh8Cp4/1z/TylSLWRJSMwgVNfxCNUhavpea3nV0sJ
UHsEWUfOxZDVaBMz7Yqjs22lYPOwffanGEz9NzdxJpSsxu1ODbiQTMsdJ1ejYpywlugnaXecfIdy
+bG8oXo8ygwhKouSptQDTzPeJLKSi8/J+zy7vRMAqA1vpdBmwkH+b9dqXoRPzujPAGkUCOWxKr83
dw2Gs/HJkrWQ9ujVtGhhFfj//k2ZnlK7lmah5FgbNMQ5+q3LfdSpxCSbf4z5T+0OU53dezoCDoi9
MBryB7a/s8GEUZLyCzC1D6k/gMoS2h5TPW0s3ugZedG87kBLgg1IasvoGyn+kVSJ+RGzzNy+AkOu
0QQCm5lUYQAkMy354LUkAVFqJjd6wcCPFauS48SKUzLx/tQ5OTvHiJAZ7q5lotsIqJ820JbtT7G3
7462r9vKavlB3n+brVoGDhTIFsC13cfBffbLOYjZJLl1LZrUdT+a9ElSpOf/+MY6sK0Y9klIP4Dg
7CzZ2LT8aH2ef9vWHOah9+yXzZypT2Ceg12pFYU2ljA4bCDYV3ybuzvwMTkZ4Mwv+uPA7PR7VVui
2wDUu+tyWPkxS8vqamLS351iM6of6TJ7sRUdYVBDkXRLjFJ6HzlwxpDqSq9TjbwL+ApYz4PPZ7fR
J2GURHSv5fQk4+Xmh3/AznT8INh1DHz3u4IqLPeZt35DHjnpdu4yjhSZZwEu4IEDhyQmkE2G7NX1
w/h5eg/W8eL1UGnjMAzWUSnYWAFwv1pW4HiXjn1OUheEb+E4t0tpyXxncm8mxUp/jxRhkB//9cOY
1OouwpWbUuPtv+D+J59So96Ox7irCc7KgJzGCcgPfrJkt1N4sOZt82q8/D+E6xwJdtmg4njpJuj8
jV0mKk0rIX/zfwkPMAUyz7H+N8OWukJo3YaEiw1Q55HYBatcaDf8a1uB9vyInEQESnY7WsT5A3zL
IPu5KiEoULw5Ecg1BNGH8lcRZc1iE0EO2mU+n+8lAN7F7Rc73msLLG5QUZk5ODWoYgP/G+vL/i9H
klJQ8sn03HIIV6MMe2dqMuytoueW/el8Ilbq2Ns3z3O0PBf3rkol877nDVQvPjJhCHsOXOag1izo
K9zAs18Pg2Uml7YhiQUT68NyovVreNGRM1tghV3btBmPru3IsUKt7Gfe1C2NlpDxO7y3Jz2zpxgp
11XeGfxSw+O+g/H3mhGO5DadGZi5Rg2LBXMzreJ98y1BwD84J1ro/zPaaTw8HpQVocv1lRl4JzSQ
WTHy+FXbPU0b2MC+2GEiUM8aH39a/pa7eNtOeivs12YFAmB8Gxi6eCWYx7b3gC4pR2tYfmLvrOUc
XIC3+ikyC8olGDWCzYwJWo32Z35GC9tcfAsMQZ+E+sqPL0ZrT8qE0+9tcujGARECUoztu/KAtzFR
VqLBsCWc+khBNI1GIRfXgXdygxS5WA9ijTRnkCcCjZuEZBjvgKlmDJHgAg0iA5hMnRNLC0s2EAHE
2ksEZa34l2wnfpE+bQpG8YkS9DgAYCtpPhLIPsdlonS3HZTXpCxz+x2bzpG5+GIobtSPBnqvUGvh
/r3m3znH6s8oRSZkEJD4kaSlOHL4Mj67uz+cV++s5SAq3hnlSqQ8R4EvqUB0nXa9rikdTA2+rpYp
R66usLqOMUqwi8RkouUIGcmLg4gqqdcpe4ovGRp1Thr55WD+Y4jee7drUn/Z6my9qDxcCWTuzUql
Fj+c6aw140OVAfKdJtriIRMSRUzHNqEQOXOhlGiiusxw5DIAtQwlnGSly01OBWqwwCFSbx7IEEgG
9yamQ+PPtbxwNXe0j1Z3JQvXBJ5NTNL5uy7n9EcWobXC+mMFsle1Jrp8V2nZL1nDWapZdRCfKBmY
Ns0BZEK/kR1kzohvsXGs4FeQaPB7VpntNZXx6p84jeOMHE1qs/jEj4Mtrn13MMSGDqvoRMzda3cy
YpAkbLM1SJyHj+nIyf8AlYzvTSyzOM+jsIMEke7Ujv2xR5julqrTLmx2Ug7Cw/bluobcPliSPMks
Fu3Zp/t+3svP5ITDIagEGK228NB3bBj+T83MCp6OcWxPmfJiNqB7nxx3B/XTwRlHBtrr7dInNThE
lDlHft8GS0o1Dr3evp96ax1zrtr5yqiznvsEpjFFP3HBBEQGDHdnmOmJ2mtb2sQtFk2H+n2/k4me
pt/sK0dv2CQkU+zDUNOkdq5rfnh9hatEm5QC9Kww0moOj+FTV2fDOO1fsYVgFtCE1zTv/T1DR4C/
FONHeR0zzgXjAqG4xSLE5MfYqxfFdrduSenfnh+gXetCdtDyF5G2Oos4Gl5SsREGrK8Ir4619y0P
qGWHY2TDVnw1h51g8o9JQ4Vbuu/0qgfNh57ZWywQMzcP/lE4lwIEVq1Z5xkawpN8gzzFU6Ik9lOi
QLTAipgI/nuB6VjTHgeUrQMKySlKddaKIQ788tmGTj1DpvS6ifQGWb4X/li4w64uPaHDnl6haibO
C8FmGekL9wkyWwrCv7LYg5+yufYl5kLxjdmsRWc77mOSsL5Ep5miBe3UpmRtNVbACT38tw8ou6KE
H4Rtc4LUU33/X27lgHC+1/pJxk8Jd3z110AgdFszLNoVBEPR3o37zBZ8LIgLQSCMZLsaXjRm6ZYs
Xa9YnJZ3szX+++lTsbtgjwrvqON018/PRH+vGZgx40+yLZUYaZtlAvBsr17x0jSs0tVUi1N/7Hg9
2BHhbpvAtsUH/hxYZOD7oMhycuxf09lVcK1Amif4/dM6hmMJCvSEiWXCvP4i0zjDPfIIZuLxeoyd
tkvZZ/n+S5vWGvpdPZlrUm2BRPkC84afoC2e8W2GeCxZ9IcR8Sc586Fb1uktxJ7wx9VxkH/2jWRH
sD557OlpE/7JChj3/zQNg4xv0NfOsk1qnzxj3E27nVr7sMhM/F/vobc4veWjasY9zhkcnvMws+6N
By1gWyUZCttTeqwmrOxTjkbgh1c163AArRG/RYowqbMedA96WIved6YP6IjjuR8qfcv+whZeuME0
fInm1mkOq5VIqbe+gPMtXq0I9Pw3pQ9XlBAnpvju+KhzBY2iBkchvJqUw5MNLHU/y1TDLpiwgpAw
mXrEQQFQU51lj2EMoWxjijGREp9PwnPRtiCMKui9hPZCH21EuVfWD9ghtI99KcQtw/+OcG2muUBW
zeDupqBcIpQRbpL5Ab4pdvyDw/UlwpFQ3NFuhhtfC5sFqM/+m+sUw6B13mocr1ornqpwbvJdNneS
lm3WsIpusvr2u8RYrevcoy+FUQgELJZBI9GumjpaBMz4gKwDNH7B6wvwYg1NDt6tqCeLa0bAyF34
VWrlwol7EnKj8pS5mQNC7lfrt9OgukXZm8SjQQq5d713zaxY/fhLZ9h9W5xpCBi1leYoz+2bwpZD
RL3SOoOFHNmuClyzNh/15v0Zg9vjoFsNy9vlg4nTLETu5BWxqbF8ahdXJ+tIIZEb7RZ0f+17PyVE
IiD5HTNh3Ck0btnS2J1COtdf2H75UNaLSsotwkK5A6Q6X8kGgMtkLUOUiANYcC1Ry1kcJU1aemnw
8S+B8mX1MZEFE12sELDqDbCYMqBnOqECjYZYgsZuzqET4NCfTyNkTxzlxHIUae5aPYnHp4GiJShd
PHhTQUpZphPnAyY+Yp+fIWxqGgW2Wx9xpMvRnjgSS9m/JecXJNw6hGLyZIzPxgY+HhaB/YOGOExM
YqZx/5O5vEWG1C4EdEgpYRDFI/Z4U8TMDYU794EQW4RMpHi6Uz2htH2LEeoj6d3p0gDa+OiXfDLa
u9WDjHdqCzOCzyQ+sU6xYh28anmh+Wlr9qdc6btQxG5utgWqWuiV7hiY8uRU/fkfioMw8DF4O57A
2l5ExosP0p5nPZ8zQbsCa7UuKScchh+FuiEAdPvZQ4BKlj2qtVjs0KcD/4t9yexQmBiS721rf+mv
qrfAK++HWwz4oEOiltLQ3gkMFxHUqRus9wsF2MHpRPaIwfb+fTTKgb9KXpAT/WMnYjojUfj34i1r
Dese0Lxq9h9Kc88tq+z4TiKpDypMDa/5ubg2PZLwnNnzmvKHFOEZjAP3xCEOkEV5GxVeLMbntIFe
BXgXQO2jbDVNgZa8BU3OpVgemjDUGdQzIeRKNM+V0ihWkhXXIiO66V2Dt0ioCgUMvqRiufy2Clb5
fnteIFChCL6ghPWq0Jm6vkhEbJyCaSgQsSXCQvqXIXg0C4BNiMQjdiCl99ro2puoB6QqpJPTq2KO
Cox6ys796rHtWQKJbFeYiN8ctYVIye7R9n8Jv0TaqqvtMKHPBRATCPXR1SRSujrK4KDp0XEjnzHj
0VWZud+w1IEFD+V+g/vdR9wgJmKZF72PWFQUyVZoiv2jxZS8buAsEeauFcWpxeheJN2v+a7oohX8
RbGOQrHTQolfhxEUd5EfVZugyNaVUgjaWpcpObqPIh1BHKyX5WVDBc7sE6fhraM2n/TRcoPqnzHK
/7ya0eJDMpj5psUa/rqut/EIw9u8WwkTyQNN6Vf3iSb7DU3xC0rp9RiiB71w4wR+B9tK7V6CZrrn
34e4h1LY8uJloPBaq94qWZR6zIXvqIxji03tG8QFkoq3U6EWaW555/xwx2AD6amXaVtIoAavACkw
crMrrk1avGrjdrUaseXi1eaDpMFCBeV0ofIAIt3+zlQqo7wYmzzFETDq8PJBTllZH3W8htyjnXmS
Zog+yugjmapewbrC4EdehjixayB+z4dCx7HP5v/8Qt9+N9gYkrE0tQwtibhOVcMgge1ugBGqDqeT
eijTTcuntF3j3zZz9bhYaTAH4cJoxMcJWIsAtOLec1UjomwMYSLh62p8KcBcplJOE0PSYoGD7ejk
rw01hpHYfdx2v2EqehZFROTtT3A7hhHyJAbi8ldi0WDORvXwzvvSa0YqCZH9ZcBv3PHJbd59/ZRA
IXOzRUZlbtWTRCqXPXfnvqFqnWsRRYj7438e9nbaQuSdhGjBx1VYn5LqrQPYTIVLqKnhUOU9SMgm
5NHjsaOLCD3C0rgKEC2LphsF4YzjDbx2CW3b7LECFw42gVFyzivSfFlBE6YUAlHHHkTG4h3DxCFN
7P5wxGKnsU0VHhl43WBe7Kwxy3iaHBJxcyy8r3kwJoCgE3OO5q4xrkONunKjdkdyI6s0ls4PHGoE
LO0TCqW9a8ONqSF9tP4aqfopMrbSsPrOqQKZltW4P0leQHIt6VLDdCBz+6MfKMJ1+Thz2DNlmj1W
3T1+ynrYMshWQpJ/PKEjz/+7saKbPm+jsEx6ZiDQj0a2Dyywoh9mPVoMHGNcpce5r7ORxJYcxvOB
1wigP+hYXRv1Sb37RNDnyFkQRVlMOa/WtVA0I43N99seJ6ET3VCZi9A461drHCpLmVpyvgqNWncW
u43996AZL0QH4sMExA4wWkYCEhPeS0U1MApU9FkE0QTjnYk8mSWLvqLTFycMPva7qKUFk2S3TCff
tNIjg6o/+GDgfDqEkP2P3A9cmkCAc5ie2wZ/rpIJ5Ap+nMFwUXLS0QFV0qRBYGwitIAA8m0l6B3r
SMpCqX15WHws8VaQYsj5Z37qtWzZcW3ptxO49uWM52A141zHSwKt/Xr90pawvVhIywjLcqSgqg+m
8OiqR1IibLoTmqVJM6JGD+0bk6iXoVzvMOHxdz0+3NIKmuXc6Gv4JPJpvEkErXYSkyF4E/USRfDL
bakJ+l00+J9d+SsShlS22joFFe0pqz/cMc3Wt/g3bP56lAGAfOkclFg/5q0saWNKOToxlidHdmpX
aD3Re7FsoqVpMFmRBTmkE5/u3zMTiPjuzG7CF/IKo257IydpMaWDeSKUEMLF/sZptiDMthvwlt/9
ujQXXsDod1gzp6rYcZ+M3cnOmLz/Edd7O6kz7aQtfETfNEAVzhwbFxuqI8JMzMK5DsXJAT8Fa51D
yelinWRbDF/BiDC9AsAUOK640EjYb8P7xIlX7affq6jdENskifrqL38llERTCqZG0XkRxLvrPsLP
BJCiEV9BICsxGZbCD8KAjUnZeAxmX6RuABVUJnfKgp9O2gnWz6LgpvhyBT4e2QUq+mha8ChPUnS3
ShPHxIoBl22TeLto5bGfCWmy/kN1kyYN3oIgEwJ/CayD60oJVWMyFU7zEWDZ/ctVJXl73o/T13AC
P0howhONJ2GdzBZoAhFyGLpRDfWMVKZTdfl5lVDQr/tRzLMRb+A2jLjy/wyuRrzayJLZufQVeHHP
PG+U1N9cae250V52YmToF4tkJv2F/rqswRsZyMciTcSfkRV2JOEAIiKX1UqSP9qt8zxmGIeob1xv
zR6Zyjf5rmKRE4SMMza+NG9JLg0C5qX48X4gWYOs5XI6LiwubSCGK5Y49H6t6IEHIvivxu2huGgi
ET4yHar8Uh5OQb+kCUZ05Pf5hb1i2P/CI3WoVtvQ39d4i8wUUe6swRlaH5tzAWxGR90wFiBC2gBJ
73BLe4sZAcXxpOahh/dRphcrjQ0GpLBo1FdBUMc1wCNKMbx4uYI3TjSOEJHH5j3Hb664I6QoSdfc
Z0RjdVZYBlvXU60jwKN4URBJYwIE+6lAANXdNPdGbCkVsOJARidYkQMG/Da8Yq1A0dTFOlrxqUiN
HPHKDNaXl5NDgUs3W2NoKPyFeGoDcB5oxCPxCfBqfFPaaspfYHT7A0zMPOgFMheHPj3TSpTBFir8
JXs/gIXyxpdfcCh5XCNLHRlvIQVIM7w8OpSi+KhCDghEO5M20AYZlwRwl8a0kFC9F0k3Ws04b5hT
szcFu+7YC92iWJddRV20IpqgIjSOGeYtli7rEZkud++eowT6fkKtj0k4SNW7WO6w39OBsw5qogL3
6kNJwSAhETkIhCg0j3AptkTr5Woj6ASEYEET4vbl/bER322hLuZTDtJI4t1FWeGL6xTmVgIPhGgm
DoZoPVpRgZ+nlqa0Zpqbqh6RSiyofq8UBzOW45oiYaX58brfIT6foqSZeTsjc/9FaLhKynICSgCp
DNpx+ToQVZLt5hdyb/OQ2K47al8KMGY9ROSi4leX0MAby4eogqu6MhpR0Rz8O8ovK8MqdoEuVwTa
XnGhIqck3iVI/KozXMQCdtdvDKtsmXB2WQ1Vn4SWoSInkHUaJC6eDP24evlaz2OzsXzIIk4I868M
zZ2PvnOgiSJA/aa6QuaQD2p6nqaiwQFwdbxKYmMc8+6f/4dBIX5w271YDKuR/qvdcxhjWY5VrbOY
mSfSNL4D2abYhkhNjG1BslFHC9oGdnrQiGytVvsihNlKspWwv3xcT3G/mm/GW2TMrQEkDvWOs/Zc
DjgcCUObun+L5sm9Z/AcGxM48ULKKGzgjjS1lpGAzJ/j4Qy6FFCpu8BR2E1XFGMi014Mnb0ZF5mY
sfqB/YFrZnVGdfb273cK/u0KWmDUq4YTATPMMkdxFNlv3bLkY/NfBcibHOJHGBRVJhvxigthVYzo
SSWEw/RzZ3WU1oA4cPVXJr6Kwkk2qaS7+pBvIO6jGmyrtcvDwHcModw9qUfWWzN1UMDnoeuis7Uc
/jxFLG2SWCt9YB6tzOwH4dxWY0cZuNUFPSq+f88f5++YWMIX4lxBoITEveazTvyB5TqvIX3b75va
+t5/s2Q4i18HbX+lppnUzivWT2rKFE+DSJn9ihjd49QqUUZgLRuDvV1v98sj+u+Kux+VmsNil+f6
PkgL9EMjA2eAVrGbTfOoka0Er6zcWtBYZbAS4Ew0ufiZRmeOoO6BI/MFQfDyGztygdZExDGlkrpl
UjXrqmgRB3ekcVq7fh3VomtUUywltru3SlRkoaXiJg54N0keBj0Jis5N4Fs4lS2fVsMrJ3iv80t8
ioHv8HjLK/Ixir5UMQZ3G0vPeoVC+2FTv66ZKHz7sestbW15bHNouuPF6I0KnMZ9zXCT+s1WJUrq
dlB2LvTx3P/Y0DlnQS0bkr79jt6ZlhFXch4TwjjW+EwoobnHn3Trk7ff/B7j63rstbYeo8qYZ62d
tZvhWc/ZWNY37iIv/VFfICLLDrBamamHZ0+PQNGV9e4kgfLDBowvwFWcaJd9WlODM6wgrUIr9N+O
z5IZbajZXE8vY89PekVOleWRqQ7/gd2T28pr/j5e8Q0iiusEu9RdyCy3/236lc/IMiz1mRWLYi+g
aVl780z6Hm8H1ZJgbQCHYAGAlC4Ep28utTNXlLBpcl4qjmrhnffXzljRbOmD1WbVIboSNtNa1oBS
WjMWD6uU1dQEKlW7KfjnkJ8s8j/u8rJC6lV39v3MEHfDNmcCAJVgiEmLB3VfUDkfp0953Sa5okBQ
FsXwu0I7AnpkHLTE559Q1vPlHxX0xpCgnQ5/nplhTWulLD1mUDC4s/NAILiiujsYKBw2tfuOmGNC
S1t4rJ5jNxtAsPB2QLcNZ0rm1ZxTH/qQFqPBPeKuBojarDnJP4f7A0XV9IZ7m0QXPOZc3GAgOdZ/
PYfbTWU3grNaEtcoEBrQzRNrBZ7Jxg3gCkOrRWPUUnRNFhOZP6A/ENREtg4XS1yiLun/yRuwCwBY
RCZJr9jo+rKuZMIVG4LZX8D54xEEGfUADtwpc9BEZ5NLCH/feERveLkPdHyHZQtv9MHcgH0CoRGH
azdB0I1touYT4DxnJ7PrRVpsjxpPpsE+xMhoLXU1DMAdM4rxdJAHRMXnUS7f17KQAxbL6IXg3UX3
n7Vgyj1Hu7/a9t16bnXKg7akfc9dsZM8iEnbOaHTVabF3QdBq4mR8N61okJsdEahkSR56E2N7uUF
WXoHu1s3aGiC9KmlaUqUbk8GpFkL4AZuZx00ZgOEboI7O9FKY3LxIV1jje9+3vHG6jIlyosubgjk
Z9O1V6wCNrykJVSP0PMl8r1OfqBmCj3K5qi9QDqRVCOjL6FAHge9e6ZbU0dGWFkisGpurbfa5C2F
DxCazzEyRNTGo69m1qo8kfPNTa3xd4rS+G5xCpwf90kH1PZgaM2lJSY5jGX9tbErwIavsz1HbyKy
7eQ4c+aQWjz5GHCTNP6zMou6X84Cn1iGMTKM5xReo15zPfGEvf9eQdpovDLk1RfnOM49lF17uyJ1
EQKzO3qosnlY7Pr0AZAQOn4Aqe2Ul4aR427u3srbNQKxGNNV4e+U6azy6rSUu0gdE2AdNpRwuJrK
xX9n3OUlLTcQaYwb074kdPaPO6CoDjC8Ev/Yb7YziyRz+rcj7Y/Uuv81kIy+iN8G1U3x1yX+8TTO
WSRNk4+slRUEnf9MU5BSzSi9TdK6jf+qVaSsdbQ/IME5yOGhth2ZNBQrMZDnKRSg14dVFYtA1ccZ
cjS+9I5Y4qvSRjY0riXiddPPmvIMH9KyDvBdfvfYB7+r6Gs/dmCTUpDKgbDSfPO+Eo8Fv5HkUiWX
jiuIgX0j+OZdgq4R/HkYo577dmKZyRh7KvIu9qnPSv4g12gjcf9ZVsEcCMV2ulubmnLTrCt8I+nG
PIQBgIpo38d8CuwnBHS73x9eIbo2WCwAA6jIK2ymThv9qHmln5kiLDDeCOIK3qCHj01bGEPwjUYN
c4A4tdACHz8wjEreUjYXf1gQS5qVUbtp49nzAylWlFBuhe/qr9GI3t4cEzicZ7Xc1L3W1Vd1d94m
duYYew9jxkrkKRC9eAg1I+hvGabORxrDnm7r+pYeXxa0V3o7MjR0a/u6rWWwgJDYMlUbvPFPNfYh
kU9TdHeu+xbmhgCN5sKZzg6IOkmqGDsQQxkAjEtg9Yidm6JloopY+2zzdIrl1+KEvubpClthglWG
SVMc4XKhdz2FtEUiTYIjNSb+Rgupxn0rXDzOWZe6MCGOlezMYWSeRYgupCN+enDLJKq8rbVfwB6m
/OIuw34tsu1pZbpkYqjI1hOpMCcn+hWrZ0zCStpAxTybao9McWRm5rRF/POlBKWZ3VVdbUyke4sv
p5z/xUFfCbM9gvcIOMi15IMsild1xRbi08zMMg6NXnfByeVdUnxAOGC2yoFEduxBU5cd2Z9tykfl
5RqSxWU9H9OFOoWsgE/CddmztbIfbQScCHsJrt0AnnwwwQI8XdXmyelsYkaLVDHeEeNw7dD6QpeD
AOYrAmJwxMTtsyy9bPlMz2eYtgx6CxuKS6F4iFT1GKmIv0wgcdR/d3ThVSsGAojp4Lo9btZ6Z1k9
o5FeZ+dInRXne0PyY5XGbV80YWjViV4WTMDnNt1Zg5dwiOMwXWpWT3t0iFF0obnk6u0Tz+jRr4gq
yuUT6F0FNJYxLi7GgR6jCAmP5TpBhCUqeREU580F1ia+UZpWKPDDfa2golsylQX+cQ8PzCCa1FSi
6qnOZIuyA8fA60OBoy1osqk7TyYgjwCoUGUzUdohNtsh8tl1NfxajLeYmEIyjKurm+hGZg8nvSup
luAPYZewVRvq/le0Z7Is71mg46EzqsdUPy9iJw/GLMX5CiTAx86pr8DYxO9NXxBvSqoKe3MxMuN3
hYwyuWpPgNz3v+ADXa0Iq+9n4GgLpGFupz6C3MLxbDNRwRVtLQtCFe970s0jz2s2sXFus0MrZEho
9DJnMvtZy68lnAMqIIxPcAgXjd+dwzgLlHIRb3eynLOx4/sCNIldWABU8wXjdNRjJOGAhEdJ4i4I
u4se+SDukPPGJBrpajboJf++MmN3SeMk1HQ9cPZsUl4b28Pv1TYy3jVOLYLEWEAXv1yiL5NhRjOU
0Ru1xIyWESO48ZmYmHZA7vNAltP8cNTrPXC0tnaq+K4eIbf+2I6kee/zqBx6xhID/Z2VvXHNbYuL
poK0f61xFRJyyoL1YF53zpKgfMN53qvx1ilCGSFLAP76IfVxx4mI8JnV3/uu5MjqT1xA5V0vdSa1
ZmiJGJshEyOi1n4IZGCwqDzTaLstPw2mZU2JJv/0qBuoUMDdEm1V3jfBO8a9wHbHFFNMaqCb7Duv
t7FmbvERJN4HpSKljOi5CWmFWQayY/7WcB7EQUvEo0dOaO4VuDHhmvbkNA56OR7rC+yN5yKIuEyf
La5fsv6oqjF/0A0a0Fj+yGhwecmsYP349AIm/il3ah+lWTFc/iKJgSyWNzbgMSZJ8k8kEOnJ+FgB
LL/Gu1urMHt/mXppmBPayImvjqg6vm6QVRdeS2FRRV49vbHZ3L5yBurIREk9O3PBjhegrFCN1Ryo
0YX2tqmkU2he71DN/R30WON7ccN9eVs+wG+2KDcGS3GeJQZ0VkPaox9fln1kpv2YpH4pzrLcNQ+1
nJq6PZpBnIuPA/HxFvxSz/bPzuW/sPBXKMuwkLr99M5l4GHgOgnk5LoV1hCmPocqOQ/SbiHRlIaW
2oAWfn1Js1aFaAIK5sdi4ApLdzTF5YtRpNXeqysZAYSB6WX/23TamQmLM3jmXk5qtO+j4Q1mNdfb
jLm9M7bpjJA6a4ZkWT9ARWby1tcbxUkDeLr3qU4xF9jCFNuI0AgOL+YsMkG3Dp7hUccGNCaEnihm
wyPM5AjSpC3bTRnA7mqhIdz0AuRt2agL+vyKG/tElVbDdxqQp8wDM38u4f4nJ3Tn5TjHYLtzyNu3
n7ul23RgZR3krAq8Kw6FkGiQcd3YHYHZwMv/01kwFj11tw/dGrDWRM8r4p1elPKRkvbIHyTEjfzL
Y+qxzonyXl+A6M5rz1107QS0vygwXzqf8flLZRysBNK2DDwnA+7yQhJDPW5/zAqp00kqeudtAqSV
g2J9Gc4L9/N3xocwAbHVCzXk535dxi2qZU38MMyanSb/a5U8XRLtJYviLX+P0pR/wwx7sMdcyfvF
itW77D2PSkp8371g7ZIm2RYlMdreb1Exp3cQWmKQnIEtdwUyNffaOnVbbtB6paDGScnCMdhTf2O7
grjk9P2CjB4hLIGS7gBLeR2JqSKMWdJDJTazp1ndVWwTXGTcCSCGHu+XEa0ckVKH8X4bSFVrcoxq
8oDw3PLJXuTEwDmiiWrQtXljW7QnmvTMEK0qsrm2ctY2rVDVB5VbNluAxITAce4pFW8slKwQD9Wl
WeFBzwaZQXJoRMCUGuc2gbv/6HeFFpERzvD9eANjv746NDWzRuVQSsRg7/svXL1kisYXM7plWHqC
DeZ6sf4B0ud3TM31TlCGkwIgaU+fw9vvkx39i7vWNcKtQFLZl1kPhIp7HjhiQkY6B+5WEGg1/WJY
TcXGiWKgXe9961ztIpPeprqKmuP2ewvU0k8j6V3dsHVeDI19n6CozdhKczLd7JD8BEVhKpiJxp8/
E++AwCpQh7jVdJzarsuLRi+/VLt2w7fefmYD485qkQcC1FSZcUkwUMfpNUtm43Ox1VZT3+ISx5RN
DsZ1rMWCrom/90rSQkozw3/7FCvbuTUNKpGppNRPi90Nh3AXPHRMzjyUFTnJsHRwhUQNckBKqiav
FxMRDCMy73cOut0rsWJakQZisdwoJmCzro0q+7cEuixKmKyWPJmJy3gWMFCTEYNZkFEeYWTsq7xn
qZS9kKOGwbfO6LevksxOFXPUaen2s6GogPs3al2+5CCimPTeRqdnmNw0OaSanUO95k7h3I8A0hqd
gsFM57z8gCf3pgkgnFLqmY4PgcSmCqmDIdSMlTla4LYhpqH8gEsgWBgVrduXOVktOgs7rOIPml9P
85mdam+lzutDYviu0oEoZ0g8iXhFZpRToZ6R8JJIIowx2g/4m/CG39cdKSVxlp/SQ5yl4ukqvZAz
/DE39kCuoIOouopa2q+DcVWkk+pz4fTPlj7IzAAG6FDpGFql7nM6zlvLORdvTvLDgTRlj779udqk
qrdhMddfZNvbDEaEy0gvAJLLD/mZyuypL+cU+Myss9rgT4EA9fXIFUQqa1BZ9apzdT2V8Ll7uFZB
MFKaVy0hl/l6ZinP/BXoKdFlYTlhEVm4r6np6Yg6fULJGCDnHJs29FQPM0KogJs7TP9uKIM4QyG+
i79SGU+zfhhsmQC6Gi4lcmOq8VhcsahGBjrDTZ9v+cSC6hW3s3P9qRXc+5x/KYcb/ANyh/WwZWaP
xylphXMO8evBPNhuzma4ntYpvx3neitkNZRAtJZ5xX8Xn9V61+iiyFGP9ANRqoqX53faI1kWMb6n
7XrjFllPkR6KmR17TrYr+AcJttZUBHmmR40UY6uqEyzEN8HRyOLk3TgCXZ/B3CPsoFjvi4bvHpDB
qFA3QnxncLiwa723iNXa2nhRFsDPBritenc5zcnMFZi40ztMuCf2iHMeiacsC14yaLceTuLuKntK
44DxjEf+IVJLh1l5yJXfjNRtUXwe981b8hNHq9XymDhmltzCuqPJTLgsyiiUZm0PfWpS9N5JI6Rx
qKAW7x4HvmzVfjpOJcT545JdctqDzB+rMLv6HcSuwycN2tI/WjSc6M5eMYn6k2MRqQHlmyDIlYLZ
2SisajqwGDPhYRamRBjvy1MC0ZjpZx/uon6HkRxDaPjL0yfPQP13CAQGcBQ/C5ESC67EKVW4PNY2
UFmBKHI3E3EOJ39izegzKr94PaVNgisEb/udYY1ezAvEMhGONC3XQOpD9GkU8IKKQZncqojEcbeZ
AswKB67LZYgDJCR863n0LkZ6A9jQF7QdEVzMsAlXMhR6i0DUNLR3dPdAZWIXnhU//w6x8CqlWcAc
dKfyvkS/XWdf/l9uQ9eRHpfZp/NHrGlzBrt6jzzWlyT+7a26+zm0VKN0V1EjhBFPQIRLgY4WzcWY
dhXckfmfQ7prUI+8p3MWEIxcBpt7WptBUEgYZQ3LkTruPk4J0/V7nCVChW+pFCbbc0SkKJaR9JU7
IMBNL1mtLiTLIW0nmcynbO7Pjtt9Q0JE8W51YE331BHN8OmFvyh4BpiBf9yd338pbjG6cjvw8DIy
nZ4yfiygiL21JwaRh6ROZ058BYY1LHXug6erPjhd4bvAB2PspTGj57ejX+gd3wSl+CJipsWlVYYd
xnQFzE/k+bwohPImox9SS8I0LZwkkJQW+OZlFe2OBm9LDxRiQ7Kl2BAm+H/pPCukYRiNcBQ0jIuB
ExfP7Mu3KbrEtWdGlPmOyIJYtbdJ4Eg6zx5IWjRLiTrbyP4ie3BtaNjbjdMizZJwxaShvIaVHLhu
GNim6mi2PzUAknimlLzoqXQ3H6k+3kfcncikRem/ReVYapFHlfHcG6IOik9RJqbt2k4s7NIV6glZ
KOCEhAopmmcuKbZ9gHqxGvtOvoxdG0/uWlUhavE5Hmvo7FrAdNxgY5vy48WZtkxOeMnng2yoyQKX
JxYIdjRvOLUqEOz7csVWUrjWWqga6Gbiyf4GUa9uC0Dvnt3LjGloU5ocVgDRxJgu7iOfoB50RzbW
h2qCZ3AWegNPCoPyswxfquLUj0qwU7KMyW/hC9y2UWUrFYUT4di3+MupRBrJKaCVsuIdFG/uQc5d
ihOopaoHxjChNAiZqFRSyo0KalEtn9KuGJPqfoThEAgqNXobgtFQTJWHU5Nv4bQzBAimxxHVT92Y
nh07UUfY0cTZoKVwdYH0R8Q+7Px4wez7PsRzwUD2mKtySS1UP2l58QW3ENpyg1vuFVmBBPpofWqw
DZgaZaJ211A/T1wiumJSOw0p82NhyZT7/+a5mIXiEqKdaSdhwCIBWgCSe5Qk5Uo0NrP/aHe0jj7W
nmkIEN3lCZXJ6rVkfQMjPiE31dHEBUTXGdUikcryL/Ka6E8babb2xoa4n+8+gZZ0/gXcw9Oburps
nR+Awq3nQG9vZTX5AZ+f1dqXOvXi2kaZfGFjS0Lkduqmhn+Q3wbUpsV9Y5mv8ozUUOHeOL82g0s7
pVXmwTu0/rEElLARswqzRDXOBTC/fK6v9Cw7gaZViSL750+9ht65r0wWixsj57pHXINZp1sDllVl
hGE/QHduaCOG3UHcScdphQVIsEBUoZQrUc1UM5m0SC61/SrCCOeCXE2RQjyHsRv25bcTFTryFmzY
/hLznkc4fTcwl0PnnLgegfcYyO2cvFfWKeH+/XBnck/pqw7LvJywhUvozEz8uWyAaIM5DdW36sAu
BGnXHhU1Vpa+OhpmGjFXWxVLyDu0IK9iARH0EipwhyLs/4CP8GHv9K/hJZETHmQ+spuy0Rk07dfj
Ky/pNDlvZuAa68EhtPeUuitj2lx/gO5cOoJRiaSRvYG4IH3WoPfbAjBwDQ4XZiz1vX8t6vHo41gW
4QTx6hreezIrmc1mjGBaXK3gBVcJbDhdkVi0BocpEy7l0MO+SoWWCjOZZXek3UiPPR24+SPTuok5
A2uJPb32/KmirOqzO762ZrepMmCI5MBCJYYyLTkGaV8+nRWPxCQx9hsLdJOM259gdrtLti3+dVAQ
QinTqdF9xw/6aUNH33LsF4jF0lpgGWcUWohhBfdnw4GiQQtJXTyXR1j9kqN678otBmlpiaryjY5Z
PsPbt+Q9g0dOvHlcNMt5lRsj66/j1PFR03iixmSVCosK1shEg9CICv+x6sbY/YqoHagBAa1Fo4LF
lW3zo8rknTbou/X0mn8mMs2a3T0SAaYa3i2gjMaHGJfBO5kEJHnzmKYtdT8h+OvEqTm+IE2w6+au
E3Yh3lH0qYikhs4deE8RxMRzjcdTL05CNBps6YdQ5o96dEJGZ45k3l20s0YpyHaw4R2ch7Fqdl2P
YGi/4jxG3dipf0c5rN6gwdCiVFIdgpwmsZDRD4ZCEXhvFBQ5tLSXCNN8/6nGX5Aaapq8J4+QvNBF
fP/n77nAajsPiJWCFM07FwAGc1wTpaH2xf1G9oRvhhrwan0rtLJcmaj5eRFb2caBxu5VsKja591E
nvPOUhecunlUSnJq945Lj8AAH1bAWccO877qCZLf7TIPF12xG1o3gXxnFT+zHjtcl+lf02A8fzbn
3w5zh3r0CM0sxe1jpIaJAoyF4vMU9p1voQkiVm2xx74RgsD48h1bmva0LQ18wJ7cpThD//sscD4n
DczFSK+piDeNR0/dbNOL3grjpvytGVfC3FbPp63S9BuE4jwWIq3d24e8Xtoparoe5GIWJ+ZKS5ys
gXZCdIMIYXoaYMWDyzQrwkxgWCLfMUmXuHM8+9XDuoNoDFgkZQCGL4i6Fx77rAZdiKFQFVkAxUoz
ns3Rf6/mP53x0Ef1Jv0yhDC2lH0FK1jwfwqP8HhbEp9QcH/Om4Zspj1iyzhk6FhIpQlPWnLXkB3J
AzAHxTyTOiYXiGBJiC5yBL0PVy4O6vNkHjPyNkMi+0qiSF3m4A4kDE9D/MSx67B+xBBKOrlUQEPB
E+vwsTCeireNw6bkjMlkR3lMFlWbIj44JlRRTieR8T4I3IEB/3xmaKpwBDXk+Jsy3RXaaUVF5Kt6
QJzHhrth1tm3zg5qWZghvXCnGj+Pgxgum7CdczEIzhrhQHHnD/K4/4cQZAtHJdyZJW7kz2E0WYQ4
OhAdjJM0Lrc5n6VP/dswYYgpQKaVK5GzFgRZrceyj8NnqQ8Ky/6uDmtZRPFFIg5mQk05tCn6iNI8
8HtPPz2tEE1dJZFcMzykOSNWaNX+3wO3BOfWsbwxXvglXXijKjxbZQXUwdCTxyrDwShkS7bq75wm
lCLH4M9JfCj0zFkfa/R+sYBcvW1yjvIK0ztLTSM1XeUN3Nct+Py7S0kUzc35KjZtINgu/eFWoNoy
Mnk1P5akAafOHjvpUKxvMNbZrCcaYGm5Qb8x9osA4UJmvMmnK7aOrs49GJnD1wYLW611XFkZb++H
lPiolW0K6NQO4O6jbJt3fFum8hpvy9Olgrk3yBvOc+8gKUVM8Fkl0YiY+BMiLP9I/6e/qgjPhj3e
rhrxL+Nq8qHcSvUG4ce4oFzyCmgnJNnoVMF0WojJQZaPQdnWPGl2loH16thcL67poPCbgDGI6YU9
qvnJBH6/EyiB8Uzq6Ldc5ju6TBa9j1zmi7yLLvOk7+vmWC0bxC4982uXorUZicmpPLGsiMCSQu1I
nhe19G3MijZ2Af5vOLI9va+W+CUUiVwsz6GFbTa7sRYxuMqxVPGdTJLX1kdeoZGY9BHnsSsb3gMG
QtG7h6tfW+jNCyN6FyKWjTB5gIw7Go4bnwzhQ++3bZriK5oBhGU5bue8Ves8I0a7CuVz+i/8XqbK
h1zvLLNZuB0xhGLQQnixEd7CGuUJvPq4+5xnIE4L8dLdWHJsDQnynAKPeCkowfXMXWYMjdkGPEnf
8KtZ6v5XEZV2MFOIqGddTgeX3XHW0d1diYZEgfkl+Km0x7eaohralohVni3CNIedyWY0FowyoN06
SSn6bgdCUI6etiqNlFfjQ72ATkT0DlEnhCq8P9oxtYxpVfb14mlhKAQZV77XevkipB1xLD0RSSkB
c6UagmdlWi7jYwpluTvZ1CzX8XlkXn7LzRVmkEdLM0Egl3vR1FmOp/zRooVyz1/XiRMuNFVRqXnR
W3xhClTsy9pkfuRzrIjHM8PlikegQ5fUDViL6n7jvUJHzak/MvEdh+3oql726tsdLtnfGhn2pto4
rgfYg259gZxpbpZoDjwTF2+zZByKAku/utBRumMxxTC24DsvgeNlJrXFBS4foZ5WBqiVU+BrTiO7
AO63YykNGqJgFcl10hnRDq9HUq/8GoIFS5ZqAJ6DerVvZUVQHvODgDXeFs07aiNjHITntscvGTk0
q2Kx1P+PG62upxdlmMdf6XcSy+skwOxfRKeOw3AtG7xRx8VI+IigpJF1/3KfbKeZ2K1HdY1gogmb
k+nMuy0tYp3YBFY4upAqyr6OkWiDXp4b9vvCvYwgf1Katm4J1Zk7t8K9hWb2Ft52jWfPl8/86z+E
kQr+FKlcJNk0nA2vdDsjT4SMVYTHL64SliETfra4fRkzStDhM9+XKBVjXQJAeWM521nlJdnPPWoL
roBnpQLuIEx7w/Lm/IcWdii2+DKr9sWEY6G0N44uwH9ewWqpFtPN75XQzjL86gXyaBEerIiSpxht
9bwxxX8sHNFzAHGn3b1m/5/zWzyZtfPVBNaFjHslGCIChOwMGH0zoMN/htZrrs5ebd/2kFHTHxfm
v5eJDsbstEwIIDbuV+cU9k4S+gc87577HMmhBPieCufK6QVvPFGBjbKYQpz0W46/IiyxgTr9X/bH
YbEHO0cj72s7INMQo66fxiVz6pVbfiqpw+CJ0gJ3PKRiwCjXDcROKfcynoosKQIzAuOIEBWyJt7/
xWpt6Vefd6oxvHfuOrmuy7nBw/iMq8hSswwT0g6cumm0yzhjVwr4unBS1sQER6wa+es0mtsNSA6E
sBEWYLtJsD9yUR83ugpTncIjyMclsWMC6vfcnIcjqbMAWcuSNMt2+sB8ZtfZUFinMPQWnKpkTzZC
Kh5h2eC7FRLIvx4qCK177I6nYwFMcEHr+jG1AoSI5aDkA+ED674TMHW4IfEEHv3J3/xf7OKp1c/5
aVTe6rtNdy78HPOhQRgjRTWAkl62UKC/K9QLs2DUVj6mIxKdGo86Uh/zuHGzDYiq1ShfY3sdjrp7
5F7/z8izVDedH4Uvzn6lXxKVrIYgHz+IGYjOmcPV3dPfpsuSwSRMnO42ewWiRrXYiV86OuG8Q3k/
oeqO6IFqKPPkYdHkA6/QW5yYqBtujFf5tmPE9kVX5E2Y/fuOc+Kt+G2Yceeq/YL0pFTOPFt6oN81
sbQ1s9+Vt9PyUKAO3BDKmVcwcObaCZxaKfSvD3dlu6YNMkFwA4tj36dqKnfrcvtDpqisXt0FNq8E
xGmypTPjQ9Dm4igMhdAJHvbh4CrXFVhgWNZbucZYF+o5fdwzKV8frsdnXIGBjpyltBZx6ex5jBH3
yMGUTYofbnHm1KykrZsfmLJ7Q27ZKGvwcoUYRcp1q/53VXMlYQf+WuRgK8q+yN5Di5QzSWsxSXFt
HPWgHEsdAuJSJrgh/km3ctgqK+L3K+BnQGFmAW7Hh/kZVOzjFjZif8NGnrSzzCEb4DNZKnvQLAHq
pF33+Nb0iGe2Ku5JPifZ8MjcK+Pk9OwAI4SA7meET/jmwx1QH5MnM7KAqm1ngDHKp7Ek2rJATk5C
cmxCXyAJkpvIi7NxqOh7RjoyWL6A5CTV64swvO3QcUuXr36eRgh4SXe57C/T/9gvI06bgh6ISxxx
JCFGmVDqSVFzhEzTIRC2IIHUY/mP/7Eg8+l4baB+cmOQwG0JoQpl6LBswtsgnY6ks9skfvKWZWJ1
EV7EaaRKzE/EfcHjunrYATGkAgQQOpjIWutk2qS/6X/Mljcj1Gvla32IlxGTh8SDkTG3gVOS25ia
+qQnexpeTQYMW2qomg3aNPopVXBGlsUCjFSa8aXYLMWwUxJsL3U5YKPsi5dRUjk/3X1C8pltToAp
N7fa7eeLZgjepafd7mrMd/kz7Ez6aT9Kr/nrXLAs6pkC7C/C3b84ol55ndPAEF3WBXG/5Kz4K8j6
Mh/9FWjsOPzMMGLb+SCfYhaQfNO3kftTLQxo0YQZzKlvbQ2JPLT3O54cA1HKo+lFC0nvMs4DfrCZ
DjRlK+rhHHWra8Fus9EFsmBFctxbowAvt+1QSNEhZoLChYPXBsICx3Vh9n7vF64H9SrJ8iQeJmwC
V/kDgBUCXLbMiYPka1U4S4HBycPewihW4K94WbIRUGk8TWa4HNowvXEIcqlArzCGvTafGPmaCLIe
EK5kMcXjKmzODfEPJ/PvFzD8vWRMAg2acbxiJoWgY9V7JMNI7PflpET8QT9wpeqp20IS7JHgwVwR
hLnicqlvzzW7iVcJyOalbMWoeP+OaKKgNRy8yIy926YBBLXcs//sz7SBH+duOTxOtP8+CyF7brQw
48hEVxyBe4DPc3ar1UReOCTCJQ0QtYYjr6hklKvE1MF2SAEjeJw+Uqzhd30OJZGy1bywXjTx/eRb
sNlI+FKyviBjlysyQgvIXNL3SDfuPIn5Zb6mgqmB02RqpPQNENeLLtkJr2XR+51IQRHJu7yKazjT
foj3zEr6Y7LkhZ0d+AyPsiZYPmmis+gYI4mMzLLJbLWh3dwyHZ7C1fNU7z4N67WJRGfyLHLS+X8d
5weVUll72CwRTPwZ6AxnkZWrPxaojJluPEP/B8Ys1KIqIS7mDUyBYxDnom0xYb/c8JMOLTSbWUfn
j82cevImjWQDodyhw9oVQ5f6K192b6DyLOGr6kYkus+VqiQ09ZU5GWAiUFka+MzGB5pwbB5QC8i/
AW/GN+yq4kNOgRjbCtWuOXGuCK7Snfu1SHZvM0V+HtwTxyBxURZWJfO2KtUkp+G+ElMu1ER402/4
mbm9TTGlDehuMLaKxX9T+iKfJ7IDmDlLXI7ErhIgeGBsH3cU62O5hzWFq5LbKWfGUGQu6WZxTYPD
39zl2UXl3kMg9YMCaG58O8WQPgtwI3S8j94nBiSAmBfBkwaupdSPD45UIxfEmzwLlzgQBYVA0eW2
PDgLZkRMZ+9juClg6O1+K6ieaEJ6PtvSVi4lxqWBRMMusG/AqjXxQo0R+Ai8M+bjbcfMGWyKg9Nc
XLUsfHBeR+Uw+uS1LOke1BU8S4RFvYzDmYMdM2kANaFVNsMRpTdFwXTkPVn1KnkklFlEQ9YLFdeq
m9pc+5q/c0/kkCa7eetbJz56/jPltZJ/Ndzxd+q7BdDKAS65FE0kVHD8AcpYrb2/GNFgnyKjAIUD
RugXv+FAFONWlj+D7vXJC0s08tTeUkGXnbocypF46D119lZ/X3GqANiJQUp+CKBo5QtzOTi7BWuT
gz7LyjcG602geLiYQM3A53IhdBhtsyZ8mlWkxUci908A/ehX+H4fJz1ufBDhuW/yWpx1wNJnGHiP
6OOcgtMVbereBPkZSijskb0RQoBoB2izb3zz/N0uv4bLQjT1UUWbmXTWoPkuhHG9N3YKtE1svy6P
kyqC8nCyTFWzV1rJwVzWorPC7mlmKQMXCC7x74+KLHsAjZpJ+Zc4zO6QM/JZ37kMGpqhCkcztwye
AjmHZcGcp6hgh3sJlmtqSrl/6ZZJyryYe3LkP9IGHUy5/Cm9icLdg5wCu3uXWhhWCpPaMounB5Qi
7B6Xu+ER13yqvUpHsncUASvu5W5kDWSAOgw+SUGfHOdp4Akx9zu1MOlPCX4BvHP+cmpGkxiXVp6D
74d2NALgFIy8e8p2Xi86CYJ1synmTdVqRp7CbCRJxq2WCbwJ4gfhM1IqTDnpt9vVmLGhFy7DAqf7
r/6H1NUXoQ+Ab4qM0YSy9WAmX56p797ol8f01cqgftKg+EZC4jnEsbTxcLRvt/06FoJ8quzdlU4U
MzAWEv33NBntn5H71lJIKuZFVbmLUNYN2JBr2jQCT6BJMaJJP7fz6jhS7HUt+QX5jZgtIW110Q9L
355t9YlAk5ipBZxPu0F4VBumI16UWnZIgu4fkdXwv0ckkfyq9Rz8LHqBloIi2JRptuJoJrqmwz7T
HgMySZTE1K2548Vc48VTEjwblR9CxFhcPwyWhnD9f69jOimsGhl9kJly3icQoqElx9j5VjtWpcp5
zjJgLkPxW9XtHX1X14/SJq2rHT7QGvHfyfYl482Up3g2obViquFu3enSO7qzpnDlS2xzqmsjJhyN
lFu/12uKnKiSTWtJx3c0tD7GjivT3a/v3p0Q5JyNigYNqJ6yBtQ1JUVYsi1583PrKK/nIkrp/9h2
j05B6XHficKCn7rE1pI2RH/nfbwOJKYmEGHcMZ7Ni6Bs17aBwG2+GaOx2kGYFVLouaPoshZZINRZ
kNG0AlaWy+PmpQqb/aTnBnLCfJzN0+UtrU9z7wY5XRfKLXGvsijc20vgrw9VFaf6WWDtebjv5PFb
cGs24Buv285SlSssKTBTVSjHxm2fbg6360E0AJmHSudKiknxvJ2I5CJXlthJpsOARZ1Bvttj/ryC
rez5s0VnzzsCgpmwAGUWIr3ilPGjiRPEGnskwaWAdBZbziu0HfxN0TpsfS7rhPuEBTC3QkbnX32c
6xOozjxqlv3DWe5ucGlpxijv6GBswMWE2RENlRssgDOOM7IMO2vab2qe/u61Xnf9+ukzAZ4Ps3XK
hUDMFylkcdUFyhcXnz7pioqXciDDVR+xyBSvBJEnuRFrkTZznxHBishJB7V1ccmt4LXosh5gvGT7
l4lK0DxH6bfS2V3l8PoXAdYkL9e2xPM/FpJxQtLRN7okkJC44haqXQiPMDhcSeIi1Jvd/n/UBYZs
ZAe3IuuIZ7L5WfOXBh7ctjgHaEPiL/kNBlMTkV2Q9HFum4t8Gv0kEabiMw6z6HJp994Crt2Tsg90
3Bo/ZLHHfrokzwaes2CU9zqL0J/JzSHq0Cbfg7RFmPpPtAYlk2edT8uLbTkLssSpQGIFJFfTzIqZ
rWVhMdLO7R7M86XChxsKL6YTD15NHO/U5EYTeVR7ddjtWPFWXFqeMm8YglYghlCFNVC0XLz45Mot
NVN3uQ7tQzCj6AXer4GOvZArCrRS2aEU7opgKZNQH7fW29yjyW1kWoHTIlHz9p9vxhcWJ4umal74
GYgpHq3KGAL0pDKeJ0eCdCFC4XG61laCWfDfjXIsLkXQafywfAZdA5RRPrvWWv5bGS7O+34N+iAj
m/MJDijVgBZwGt1o3YBuXyWSNg5+ofP7Pf7pETBuktfQk992/DUUPZLAEs0beqlN/Ohj1jDwgYNf
aUKrxixaC20ZBjdMEL9GBcT/P/4lCC75fMxVld/a2PTMfJAD21EP227IHndXOZaL1YW0cKe59s67
xmqhDd6wsUeXs8mJS2TOMwgqh/isQ9QyNzEww1w+ufFH9Y9ffb4FuacUNvZSRYCWh7ofBbb2uZN3
aeHQjyrmhS8jCP6GOtZ8D1k4Ip+JtVqKvJf8Fmd/xx4EGRih169ClA/eZYBBM+Qo4BHMbcVJeKPG
l7f/XpVdpXCKCUoTH67s+cGUw9lfnQLuDgD0ktnHlt303m2zOfHTUzjw3aoNo/CxjgZSrljTf3LW
CHMjdUZXByrdQRwLQTRD8e220ei80Y8+UfTU6TgApDCV2TmTx78Zh9eXYeUWkYzufC2V+GCpH6rk
1tDnUaUg04hEzCmevx5fCeaWaaS8QPSRILTGURnNKY/A/bS5I66YOJwD/HoWBNTKoe4JP6g2fGzH
a+OcWOH0qZLPXQ5PMcPzbMdGmGaT9EPA1CC5ZiQkb1w/L8DJtOBAYx5lgSXJu8xeBkvc3HZLXLnY
RdtGoEylcsE0BwevqTmO3ri3wgq3VVXWtOGK2+M36EoNpNhRM7kJAkeAr7XClDSyZe49h8FtOOkI
T4jiKRf/DMwfMlw9GJcCa7/6gBimBVny1EsB9iiEarwHR8cUx64CtAbE3SUUlWSjHZ+VVErHxNMp
whM7jDWfDrbcY5nJTxEC9QlwJFkG1piznERSVm+o/LOHRhFoNHW1IBWmfAb8tiWDvJeZulNTqxBP
Uh7YGPa8oIuGM2S7yddDMsGTq4T1Sf7OZnOiPlOlU1hPwUjHtSDdiq6e3KO/eDLD6e8Prtfc0NT6
4ilDrgcR5cyF+bEZH/M4qlu5xAa2Iwo7K9xk6XWvC0Pz7eNVzSC6JgASQZeJ4OtTGWcwqEuHNim9
nuF7xyXxsGpWGita2nLtCJtRS9gVV2O9qOYrRjl+Gwb3W7U+vM+6wAAlmifVuxv6NcrVDRfctjIU
wBtIEUI/ee+fBAhg+8sAzZEw1JTSt9VJ3BHgSQIwncVyiCgf+f2R+Qq+LpVnbMNeOHdgnYCiXxNw
D32ZhmPQbnOCzkaCv+DB0r5PTYzCSO9xK04xhm1qySzge2nF0b+5TRks2EYve5KEQ0iwnjOaueqG
d2qD99c4+nR7BEs7eXrsdtjnnLD4soA4R0F8o/RZwNSYe/9NgSjA7cZnBDyaMm+YpxiyFa7hd1BY
nYbDV6urTt3BtkMf+eWw72tHSb2Z8Ikq3vQ3tO9nuF6p8HTXyZYmOp6n0M3cHGG5ucveKjDNKWRh
wwmhW7KRA5mkXEc+uiceOKkQIOUSpm2jc2jpUmTaVgDqddIL1CucytJZHD4hfJQ32V1Xghli+S2m
xGZHPHrQ6TUzHZA5aQ2tkgPH1HD0E6uw+FyJATZvVX6uzMS5lC8jfVgdvdWSm/l66iMmSuJZZASQ
/TnDzPR2EoSxILP5sj/AMz5SHjSwIpHIFugiyEP1QBpU9b6riADJ0DHVuIqARgBKS8rBCbrglWeb
vh8O3FeYcRQH84teMg2uA9Dtkk2kr77TcfQOehEJhoENNJG2OqzT7dPwhY94/1TJHc/dyULbjYWL
kS8eU3daQoGiwgz5j5pSCh67HepqNo17MTUAwRrvvwMwdI/b16VoMjAB8OEhbV3wF9xIxUKkw07m
NuRDo7eQof9dEIs8vzp3jmD5ZjXfhgpjvlUF57tRxpvVxx4s/cmmoKY85KZcOBKBQjd4D/6ypHZJ
++h41aN32PHRbrRBL3vKORQcjIUquQBrrhV7mYy8NT0o8Op7LKv4LCCE4Zn2JO3l/FBIC6ttGmWe
8r1lz6RgSqdEQQia8EAKPvAmK6huxLK9CZb1Uq4xMTLoOLQgPYCF2gEItQLopDPqeidnoAKNZ4Li
3Z3H4bDQTd4JsJiJgxNvajGlFSZ6qEGZNwzvo4l7is3gM9qwX0jmd3IlTppnh1YEoAeDPgjohfpy
UnSWxOd45bLF0miBqHWQDNxqzZH6Q8M96GEwid8wXfP9kOw52XKvE2cH8q3P0O0RozGl2GBL/I7g
rEQA21VttBimPqOyCrdvBb0ME+e+RwaEMnOu3n8O0sRfCz4h6KbOs41la15KUCqsPQZxWEEDlW42
3JkAd8DDhbejyzWjlVpsnSkont06okHdC74JB0ObYOV9xl5IL5YNyvLtHmBkiZ/Ga41v2D3HR4Mz
shzsB+d6IyQOtqocI82tcvKb95u/SSj5v6IEd97vPqzWrSsPylNx7jKIhVfXqkNKY0YJZTgdHJHD
JszX9X6sSZuiqLpqXrK88eNbzs1tBLhvkT4agHB1Hx0hjR0soQqMHNnqGL85gJhge+X3wBdMTSu+
jiFphmCp7ogucHo4BTJzw9KaQqZz0EeLuvSRFFiaYsHRKHx1hXGjbQ/Y64zbNCBLKGlzDP80HfHd
nwcYn5B3Jpu6UkieQ8kWZTUCNL3SG8uUD3IdBGJZhmrRcfL/sM/mr/GS4qW5w82AmHMl7mkQR2+x
XUMT/ej9OEg0KYxx2jaW6fov54UWzhOmQWx9yQEEet7T92ZcUybLib37eRqV0575uUAXohpO849D
gA10xveQe/Qzq7uet9CCxi1hIPh+5WB5CFOJIO1m375kHL0x7aBoNoJIhOB3ut4DiER4xmQcibIV
d007V+QVQraFvZR7dz0ubLqWL4jN/LsQ6/pHP9zbUftG4KQP+jd22snrUREgqpENtIUaXZKZAC/n
u72CH67sdblXb8NPIFqaSGkn/QIIuj/kKxL6lIa/18WbQFXobXEMjIUa7iw1rhHTxUYw/1xXI47U
+VyPAzLkZWV9rcGzoziF6pcz6Kad1IkCaZNYn5K7XAj9FgWbar1XlPGm2L/5S/dfIEqzQm/MGmWn
aoTTyUPro5rEAn/mtukNpDiS3ZuRNs9Nh6lsSp59LK9qQzpBC82j7F1lkQajoLb6Gxjti+lBWQCU
pn/iVN5bI4xwEhG8rlwfaXuIiAN7Zkye7SrAsEyFx2k0jfOuqxCafV8CsnYpOmmphscM59agPvYa
2RcOpQeApzzZ8/2DGjSYVGL3jeXLE05cQT73KWkPD7qlGHNFpKW5FF9UXBmZcAi9ed35nbo6MqMt
6gInDA1TyNF7b9/3LSG29wu23qc5UzcKaw3auvU8gthsDd5+Y2RpFozGv1AnkvbjDc/SGi+ezTd9
A4c64hz8YvnO9AT5yZDM2iW8wOleGCjgYR7mZfNQuF6USScgBch+ijNTgwLhNSfu+kfzD+Sh5JgT
3Qe2fyJZvRdHQoFbcLmGHnmIvjYtXSqqcWkbvb0vwtzbmkRX5qFb74VspC9snUawDVFrVykp4TTS
kalplQSBhCduLxwmdoz/AuMUFigdthp5dN+HruFk4clC4529o0H+rb1FNvn6xohuUh8p6yL2isd+
sNKFjl/1oxd3TdP9BO+NBJxpZy2TWrhphLLBvq8+3vzb97zz6ZLmHu9cn0OfdgL77S6rWm9/SgZC
cwbIRKVDRzi52NF04c/DMXUo6iliVP74xy0lBZ1PE1B7l/6LSkJ8e7KQGf0q5hqr7hXkaJs9Ja7X
rGu173tJE7SyeCf90uZUR3Gmgk9Plu/eGKsPIjtEpkLx2N9z+ltzQ4H4+Z6nuQdcU0CV4Otl1lPj
F+NmaRxKOB4rmfERzG1WefeL6S3lx6kIXFRg2xUIyY4e59By77/TWBkBG2dGbn8uzUWvWlT6Atan
j4Q22pD2LEEkNJiJOjrLaeZdtX57Xa7jzJf+0vtlJ6UHl+1ppAYknQ93rq4b/BPJVgsH0eseihRC
7zJj2m1NhrkppEkhoCdDQtQ4gWmQkf2T5x3XlIHKuWbsjlRgnPadWSjzr/tcaJ+wVL/0KRJuvch5
9paR92VZq9AG7FZIa2obOtp+nrRGonnr4Ay9xeI91Xdkubvy+37UgC3hbpydLrZJUG9b+2l5b+8f
RUnR5THyzvtGUHHRn1CQDiTV67tG6C2AiXnkVRvhKRc1ZaiQxLiAtjhSmakaLs8Q2k+D8OKaaxdq
7YoBQ5efwFVoafJv5pDSVX6rckxnHdK6k7XuB9XRQfxtgKH/+PLidX1Uo0hQcqvpYh08QhP5XbIm
xENcP3XP7/gWW5OvvWVueOfzlPIabbyhOhNsY0Ykayv/zw5CEx7mwh3i8pnJBX43GU2PTysw14/u
9Csyru/jd2VdxsCGFv0kd2h8MPO+8eoI2pLCKB35XS3KPkY2t/oHAM25PtNd4mtt++wSsqUbe9QN
fUq+lkZ48ddUbs6QQ1O75lCaCkewC04NIS/NBZg8IIEi0Du9WIKNt2pgBXpam2YwA+KHU4Xkl42w
n3bdSym5mok0yIHs0C9ZUbsSLfeMoiybKi8YFxdwY0U2E9VBY3csk0d8gdOO8yzSpVj4N/qmykcD
HMqLh/Y77sq9RB2g/zOdFW7Wg2wPQ4KfPIcPIs/KPt1VvnhI2A5kM0rjZ7DjkIn9MZGErXaM7IYW
XM9QOWsUlS8KLeZMP2pHCC/i+Yfu2taKc37vLbYN3o0M0K84lXX0cA9C3VN8n4pxt1q1pKjaBdc6
n9GxdUg+NFTCAYnvPsSkeXYczz4w5BIcWGaZSq/Eug9bmrtQ9oAmNum6Q+FxoP9rNbhPf9HwePQq
X7jPeslknI3+6ML0FFDURI3zOyk1lEtU5PdwXP84f8rk5x/PQaV1Sh9zpv18/gY67l2VrwDD4Iqc
xlKd/QQVzDWsOYCox0bgk2u1EeLyN+hF6TYmexS1DMkLmj9JQi1jSC+VGDqw3ismtSDg4KFoamlw
BBf+KIGuO+qORNdYTrN6UOBmj5euYGtPreREjYL5aNU5qRl6uBR7Jvz/Qv6tF3NbE8hRhK6WGyWD
etwqwgIX+hxutvlPOivIDHNYltLyKCDHI8OIbuJtsO7Ty6eHiu/Q5xRdlaGqjmGnRM1bpC1jlU6H
zzX0a8rzURpuE2NgCODc3VbxmeimAScbcqqd7vMs3W8SQZc2hsnJ6xzkNeEJ4HNLDasB1WNF5rVh
wM8bz132nkEmfPHFwoGX552cse8ZZtmo1b09aH5XeSVrvc2c2jdHkw5z9l/B54uMDEogiS29SGLd
tYjCYkpPtlfEjNPius71NoHS62uYkQSDl/bu+38s6aEEFibIY9e/cSzzE17ctG7L2cOqfWf2CF3s
u6gOr4A/ZAhXGda/VOxRzYVfeECOZAI8TAOsXVIPClDltmpXHO1yrEQ5EYoHAYs4ejrwsWt5Fa3A
pahUnBnf4CvG9GX+NJZKn5TQSF5Nks6GjX+s1jfVmETOrVZXwEDN70K3wATYTJVkm3ZXef6J6hBI
hPphRQVIFAbVixDiPQ91DW/GweDqti6ZTi6X+hcj+P8YSl9KyuWlaJk7P7kDlbJTlUd8XiGAD72r
zcV3CAal6Z9OW3TuGQ6Of1jdW8iGvakDHr3lMKtXJQ3C3wdj1tx/OWn8bVfdSpTLJsvxd9lhfuQs
kp846f/ezv+2+RlpMriErHx1XEsuSNBYjp0LWcOg8vAFa4fjXLzivHzLBIC6c23mheHVIEYc3i3n
+YyYnhOYnwuArE96p/l7A+6fjgJrG2WOPngwwbsglbVSg+FM2+lxPkriDtQv9k3krOF8hYxnO1Ft
T0FIcJ6Ex1RLbC6Zd+K1rzLNHLv7a44N6CwXvJ5btn+YFFrHFfqImh+yrBGroqW92z4rrINlNwB9
Xhnv3ZkNCn/EsI54dFDGPWuKqZPykLB1PN9weBV4XiljoYHzZaYQM5b4z1KDPqNyZCtp3Qmr/6ZY
x/+3DnD+ElDjsTioo69WV23yvVnZjORdu6fXd2RCoT6r48XgoWGvoM1CaYFk52xcFwFkKAhQDQpF
gMhwPCwqGX61eI494y4Q6oU6vKdDgWHiEUxabqISlsv+mswaCUl7Np9ZF4qMky3i5oJf5k3LTO01
1oa3iWYBePI30AlVf/IwG2HLuhXsjz4NpWT2ahMHc2pZ8nb5HiW1OLYYyzPke5MIP4+hFzllAujC
Gkb3eVF0wdEQo9ipunvcq2U1xAc2VEkEzqnOGqh57vOLBPNlK5981nvPz55aFjxwPQiNIu7+W6jc
0sgzpbwDLVDVMCWx2TS2PJumBWm07FlGsmvw4kA1F8iNund9J542u5VL4Ch4m7gkvrZ78NUy3yh+
iwoDJ/I8VwAmciuyTpsHOLolpUr3BdEpk9rdy/vFCzpuE1Znz+C9qmZuJzdgc/V7X2g03/QHbB77
oVo1pKfKPB8b/hCZZltPskVqojbwTpJgOEdTZ25trQsaJs5dTaf0VHTM7XeFXqiuEHOjHBGyhftR
Msm2YRlBYWctcZLxvpAx590D6TdkDvZlsLaU1/kHlsCkmBhNgbs8BePqLXZ09FubjLfNa5X9zm9T
YwYryGO+XZp2LEotNFgo1GdQGCWl0wLa4HCjmgPHGOw6YkQ0vUR4XFaP9tNzAyRx69k3e9wn19iq
IYl1m/vq5YKCCHQwQ/zbb9LUb2VN0u8Le5SsA4SvUzfcfoPPYxIvJBtEJrg5nq6V+8i4CEGdXTIB
8TlRH2uQnKiDHHIdxVywd5SfiPc8W/3SVcDZqE1j0gtv9HeMaa7I674ErrKV9wKU1GogFWPkcZjX
Uf3jQhyhUPwteiwjDa9nKh4kNvZzq+jXhhwJzi5DYrswV5IFa/yfZg8zR9IkJbJ5NrJqkLAaonKY
omQIWNiHnUZdP54Ecag9cI2MAMPhH1GzYOyGp5YAztKlX3StFNBTpbqjX08dcnxAGS32f+SUX5ml
BjgHS3r/yQOyX5V8//L/XNHy6Mp1IqRbP549sZKRq+Ol7U+Ys/H4qxLHt2ODxNz09tDvPMxdBcfq
h//evCOOEaWGq9VWRT3kNKB6NIlP8H8gviHJHuHwiL+7gz5mNZNVh8WE0zojguR5HOMlHDfOtPEK
lXIG+60j56Y7vLJCsNDkQuzQYW4F/dvd6b0xbgcgtgFilJWNpqLF/VwLYCMK4aMpVAEkYRsQtP/i
Wqql2aTXSRcOWpBY2RMOpMaBEyF7XguyeVVIoWYn2hugfohABkn4p6lhP3pd5ujjFFa1xbE6Jwnm
2bBWZ4KL773ajZDNoqFgHofMyfJ8UqL/L05lQsu2S3v+fjBmqJ4aORO3KGk3hOVcJhHizrB8RQkt
9KgbAZTpQeM/u/jnR2AQLjptyEQ8WUij95Of1EjcW5BYS43droVqcp7mNUh+Rjpeq/y0X5iznd7z
SWghGMOULi773spJCy8QGSe7o6lMo78gFtqnv8+TlK9DjmNlyOahaR92XfKLXixwUbQHBkh0jyKW
lt1BaN7I41yqQ7grO/laP8LOPXUZaKX38lqUjR1Ol+TrgVyjp/jQQ2jLZfrrCU6mFaNCNUM/IRtu
4J8KZU07+XMzJfqWjCHr4j8/v+mS26hDP14kZeLtPVAmwPbeTUu4yeYaagsf8Nz/gdaH//S08Vmd
n8qTN//3dPJvAk/P8gjDTBa5o1ckOFH2fpuPhS3HxPQdtiaiiX7OH+GVCkBIItvahu5mNN5Do0ph
WMcHGQlQoREpi4a7M470JuH3NcKIWlEvatXHhXphLxCL0Z9CNfzQ+ZiAGbBwZFpDDQY2rOY5w0OX
7Sy6GUr1B5bRp1uyZEDi07WanuPXG+GWKMQut/biO9pcg571OnABZms2LDyRujEvpr4aJjQCogKN
VanVnLXoZX+HdcqD+6I0RJvYgtK8xDthX0NI+yQn2I5vyxIU4X+x3bxiCju+WGX2fCgR8drmC43J
6tU7QvkmLuIds+hXil1GVqoS9wodFFBl85kcZxc2BPrTspzrDdj/f7hrcp2FO1fDuWbLabxBch5O
GexwMlTHhYtzHSrBlFDbwwvcpOb3PUl54W0ZKlmgd2PIq6mtNgTRyzp77Hg3rt8/fXZjxZaZfyjc
Z6nankwIqyaYbCNp+5PXzIoRiw/6CQtzccARLcZRSP91SqQhjz1QYEW02yK71XaBXitOy5sEVv1H
3llEX3KImQm9PmHXR/sAPNyAldG1SPrAJPAjRf+dBH5xGceHvFdjz9QoAPlqsC6PhNTnI4KCfTgg
Guqv1E1IAzPoIn3hLgDMX3y4Ls+7jtILfUrLIJp7WK5Iq8kZAsJ7rwY7znQB20HruYxMjz1TyR4L
gevAhPWhdoblo8LWkbf3cBw/CBebBZ6JQby0hk1g+baU+HzDWM9R4N5UGm/n/Hw0hwzv5WSMaKfb
MiK6uTVXdZHKxy6IbmRkh0Bu3ALnDmGaaB3oovErI+j+mjbnjcxdMQAjJs+zKE8Fa2L2nHgugDfp
aPU0EIo9cOPQNq+iN/R19f7+6LwL/a+1i8law//QhkGFjCnB5JLTlQf2O2MeIETJAhb1c/gKO4FA
AZ9+IAp0UjuYsS+6hIC0cTjoPPHR+18pKrkgw5mlvYZmwMWcSd6kfFhlN1hem88reC0aCviqo6C2
uMhMSy6v39Zz+5sddM6GAmsAWV5Al/YbT8UN8s/AUiSQjZS8b7ApwQQ2XA1M4hxQczufZ50pxsYS
vBUIabMLoZ7ev3pUfEiylhCp47ni5XKjoYo3Az7/hk3HuELzeY1kDVCazgJRsf0MNgvN3MUQuOHJ
2gUrhioq7lMYJwaXe4z7zkV2idNxlJXY5kbUWy9bVhioTdQhUBDde+Jqtj3llY/1lIAHzz8MMOfT
VqYSx6sO4PBQbXUFLe3yjQCtirK5xSuVqoG7la+7lpCQcwO81zFyx4IjxsbEcAhuL44xW2QDd2Ry
LFgvC8KY3GBmzj9YzkfCKRcqV6gt9eAN07r2l3/0sV1HwKWZn4g3milgRovYbW7+owqHoapilrzy
KTAupuPiYvBQU/zRhFcoAJVqCfTU7YHJoyZEUugatcPkpsSjlmk+uZtHu7RsubE8sdZz4dyenXbY
o89e17JXhLfTqV3ag1arvMg7MJKNLmx6c3HgyTiFdW74ffKvdOgZerd9VHKQP4zI0XZql2oI3a0g
hJFow5jLFsp+2UrJ3ES4fHyRK3DNcaO+/JpXb50/jtZnsH6cMJ+G/Gq9avifqL8j/JGt5diBSyGg
yaysyYva/MP3qg43aTffiSBF5+yz6OuR8MlUFoCnd+9KnS5vlpC6KMqKQpF+fLBaOeL2IxiOa1Fl
9Y781f14KpTxs4+yPJt2AEmb/oSDB6BNZjAQCjh8eWxIFUJY04W2x8BsZdYhJgJRXEcWgvU0S0xU
u2OyIEYyZOFOW9bOfEEGJgqcJf7RkfIKXECa8KYeYJQ6Hjv6t8QIqUOht+x5Azj454jpUYbdZAn+
zJg2GWMF70MEXwuqs+naFmtzJqdKcamzsXsDJqG2FLuU70/lneATz1F0wjsa/33UnKaVs24z5eDE
SDSUUgGFWzc5ZF6UZbK/L2zgxnymtJgdvf7r6dgoQI7KjcQpC+8c/3Osc7sLhnF6pOAdjX+x8WAc
dabaWh0LSoNEtaUzw4z8wMaklX1Hm8WO9AjCrxqzvNXAslN/3L+kNioO9AwfMDIN3ylGQ35glhY1
CgeGGfUqRd0VPL9MmR9XaMeklt52w9qYkYhU32xWXBkwHhNReqOnnNnMoV0LLC/pliPoAxvYALdg
6j3ZsA+HOHMBsCa/ZIvDFxestfduHyIPRoQL8IuNO+9M37w3dD3m2KYoFS4Oziyk4p6jP4DDVDYX
oRAoVkcmUBLGvdvqsK9gXTFyPcMt+u30c6brApozihBXwRzdBA/SD4NkfCc5belIUSngCaGwqkJT
Sp3Pic9t0hUJWnpDVos8GTucgcTDTnHaKnCym+onnjOBeOVs2pF3EJ7r0i1r4SxdNcrpNHNO4x+K
CCSbzG1yPzqbtLPxuMuEyXCqEyL59Y+zKHVXnJfmy0e2ySEexcoV1QGc+di12xVxT24EW3Bn/y09
oJy+JrGM4Vwxa9KmWV2RBEqXj8JelYS4QdGVd5Db3kfIWw0ao4aTc/V9t7+ARwYQmoiLKOD2vsaD
St1qhoCKB57e1x9J8JvzwVGa3A2pffEPGrgCWTXXjn5J0BZaUldXI4XK30QR2dopUVQMwnO3+kEo
dJKlNm89FRlIsSQ7N0cRepYwJk+qmDX145TmZ6zN/MhRIaMccVzWCfbhGLT/H0AbwcW0sVLf7mc3
6l3BZzJGfynVue0pqtQIF4P7ZUza2eQyWUMXpCCFFNS9TeQKax4MVD43jFvBW104PtrNHrfNallB
WJzPbT9nt7BGdOZx8glFrbVhZX3zg4BXGjxTpkW3YKM53wplkAcloHQ44HwnuQLombKcE6oYZVCs
0XLLjNQeaAH3cnHS6r/9bYa7Jj2W2B9/ASNaRC0trRFvtrF3Cv13CQTRJbRdXr5qX3i3AKz5+XLr
A2zWe3KEgp6TK/YSEsDxVVBcEQCCsZAVvSeD/+Wl7s1XDLt1iRYmPtbHuMbT6GxyU5Zewe34V1rK
qJt6nG3kgGEoEIitky9ONYQ6jaQ6dGEgckm2QNNNhtohA6K2KbaoLlSDbxrOg2aJOkeIg26F7ZOq
FTextNPf3IkFTAl2yQKoTOFW+hVB+Md6Z1Dx/91PwS4aq1B7UuOjzMVqSOSkLykXTaD5HwiGoybI
M+WfewY71yhx7LHA5ESKDWMBtdDCVkA8+zuyjDKOTsP2h0trAW80TmoJkjrrs0P7A7fjYB0JWy8z
rrz8JYbOrIVh6erPaHdewZHc7XtN99EPm5V5iJOpB81k7ocB03jjY+x+lQ9nD0DC4+7IAlSzOJz9
YhIKY92R/gufdh4IBt7Kw3VrFv2j1KRM5GD61CAqSIy4L8XZQZRHqtRzrQnshfcn3L2GECyGNMaj
Kdc/On0ZzRC2uq8gkUq6Y36amUV9005ASUT8glFrewBRLicM6gtn6BVKXqhPQDxILxy0fh7RnMbm
8xPv9gqJ4eVXwQk6DIp+qRFxrKCf+2P21WRRF87FjN+dn9E4O5ZPaFAXZobafxkBudeiflrqzCPh
aHFGKgWV+AZ0GDMik/x/Q7A1ROfSJzeU7YE+JCvKCJRRW2WVqjlR19EL0gZiRwnAlZleH0sbesdQ
jzz6PIdO3h5ZXTORXCE3luupz6R+FAWcHJr//qMC7b8TEcURRituJyXv0WXve63d31LgK10/jLpc
1mq3Qk2mgBFwSOSFpoy3PLBR6KPv3dCOS0oBtEc7oaITskfO+6Iy/8Oj3thpIeEt7e1ot/E0PYOM
ee/Aj4e5+6mIMa1PpIKw6ruDSdUyXBK1TefRboHfY9H/36WPcmlcDTr5BVeS+F0ofs8eS88fqDhO
wnJfv1a3c8o+9fMK9b6fwYH4uSA0kxa1MAkYiQv+QWw5RMF1P7TS9DhZPnjCB+nljyDwbWZ7EiKN
6FkVi0M0TknG0/CQtCO0PjOqgHHLxmjVDw7FT7jgUzPFMdxdInL3PYJoDhAhAZbvcaqBHBYvkxuM
WfOVK2qmjUSlvf+pVbLVmYEark8wdC+0c8eKqZlIYCNJ3SdofW1Fex4k58QmCCM8fAu572Iupkyf
rAvEkTYi+F9vxPsdfcWyjBOUW+//45K1XEwKJxMmICPV5SAH+A56ozn2GhR1+t8t61Nu82pPoEdH
fzMmFLZuCOCZQzR9DJ9y7gsX2gH2ZVmlkEwfJ65KYFavj3FOZzgOs/ROpbJn06Lpd52y3GBq3zFM
w8PFmBEY/d78oL5QSKLlevl5Kelyx3lm3/3RRAX3s3QRObZlhJpLwRT00bpkSb2q2rjomvjQqVqy
PXecSGPN79rHtBz85I5tBALtXgKR9E2rDjeXijAhUZA7fCNoObC/1Td9XF5BfIwP/qzQQ1QsZMjL
+88aRbC3ChdrttHIUVe0vyUo7SkwbY5g5s2MRc3OrnicKVQI0mwQjnbkF8NbHKq67pmG5MPTQWU0
t16iywGGpuCQpgJSSLmCMUXiKKi4RVSMM8XpS002Ulm/8LbWYtL1TplwUDiq1yjs4j0ENL7IRxNS
exBSieIMtHuZvl13Rdqbdueqii1X9ZSpXQY8YqehTYZNyxOqgcee8m+oPO/ddEcel5aPd9CyCvcI
8HhnZHOBl841YxgOBh0voxkH63qWwhaneknR8xx5T46pqWIHFM1ZaltrN/YoyFUP+Y3ShV7JLXEj
vYUp4Lx4rxt76FNkKgw2jC891KZKToLYqpMEbMZU/bWkIav1GHoeXlFtN/yHWUCibGvueQfygLgJ
70kjEAbJIWikYcH58EoE0cMeP25ufUipBYJ6pgPzs0cGAUA0fwxxAGXbuxu4EbuBLwgPx2OCQubY
Gohf8uVjGsnFHJBbGONEEdTvxdvAWi0PzDf42X73giRJqGBROzOi+cYkVFmFwhEFXIFrwo/JkLhc
Elwiqz/YxfpeuFYarxgAOqtlST6X61TM5itjxaWWK7RZ+juhsIoM0YTht0bopy6hbrCmoiUjI8gQ
erHafwEGN8R+v65C4/aW4x4IhcH+4cb/vPm7glXtTHta+zMaJv2FxiwYliu9+SJcI3o4KXGKlWeS
yY8n7zwrarVldq4w0JeiUW0D9xhT3p+zyIc/qMeDJcdYM1eOaFw1ROd/LSDsvZshhfl6IegFOAwa
j4Q7E7r6Nix7qR8P8y81ZDXbOpoUiGm6ILYhCx6DNpqznkFyJXXRu/hKmXovtRQdGNX0H/kLbph5
Td/JwoOXYpQ7Rd9oge+O9Z4FplJisUp6S5h1VO6Cq0o+F2XAIVdhTgWP9s99F/O3hheE9IeyIc3K
bDse9vML+Dnar+UTSJzAE3K/c/ST8y3dDJfKa71Y1x0dD3cJgofzcR7Sa9RPWVJ8KSjXapSgf1Cs
Vebj6uqE/X5a1pQP+8pfUyOjZhtf7ypI5sV0UBGoEs1CVfmrJs0L1tQEObUNpTMU+EglaYMVIKYj
GPcQ8YnawlEqybxEtnAnPpVxRTGF+TXhhMxaIvWR5JO0+Or8LGztI79CroTE+dcAF1gCxcGQVYvZ
CzoL8m3DS/C4wFCuPvzTNSERC+vMbsT7GSQXxxowqR3rigDpJuk68F1ub6/FIV588X9HCirGPXud
1S1v+PkaEKIonJ1phPyQ2voQ6D0wgx7PKdbE0yHOf1NKIQanDZ+9ABkkkGnD4hAcUwgvEAtUgO85
dcJzDV7pGug/Jxh8/HicpNagtjIlXFG0G1tQFZd5beLb6YKjUNdepzx3GGRr2aqwTMfVsnTlg22H
Rknqvh8ZUg9Eh/DZ92k0JR7NVYMOCfRCdZTR76xkOQL6V0qf+/KdL+f6Bi09f+w0t9oaHQClqC+p
/hgsf9rTtHeEa7SCrIW7PiSDiMMCsjc3Bd0N541DXLScA2P4Ju5+MscZ5rB12Uxz6MELhz2sbfu+
UBJRoE+ZnNrdCbQ6gzzgl6Y/wR0sB+SZx07daQhp2PScXJkGGFt2rPqSkuzk93HKVGr/wlYAGXDW
720RAzVyKA3QiZdH8Y5amJ715pk/8zeecsCg/valUXwTVFD6Vb1CB+X9EKvNActZl1P2qUmhKy6D
TbN1aAHvDc7zsKF0upVvFGAJx4A3ROCbTfR4JHmzOuoGMgpG2m1KXdCM4rlqrvdaovW9s+99n0kH
SiQAo+xcMRA1H4j/PwW5vszgw3wxN+DIUcZZ54SIk/D9biX3cN1F33Z1dd25yv4ar3cQPOp3hADX
zlMorwaSdEejCCKCsfngbAro8b12LgDD1oWLEg+vUmGrw998SvX046/xDC25Rh87bgc5HTb7y/oX
BzFHGap/2Jp7E/sndxy0OF0UY8W+7P25Uv1MWLNFThassM/8ybZttRnU8VlIA1fZdynyvcOqHQMJ
EOVDN19s4VjJPOiUelrxxvph7wn7xF9fiQdyGVYvj1E4SEHXrA7/pUDlyl8UOjPigAJfh/Sv5A5U
jqpEb4mKrXiXd1ChlZyrF/bq/Qag7j+0aa+PvrlUqOfB4CeKyBbFeNR1ImORSSPUDXiFfwiRgR4L
tNBmrVBnrF6+BX/g+kOYoYWRL62pt2m4MBZlOArIWj/+L4Fc+vdg97UwwiXjjwjW8tOtpTF/Nv/g
HGLBauyUH1I6uz2Nk+91mR11tBvvaT9W0iLB1nfyeInSAYTdLQh01KuU87UDozORw2HFMmBFtU2E
R9Lx/EySF3SUwltr5C31NkfKeVGk1Bdc4+t7LCVIwJpOM4qkyIY3Dm3lGnVXeh+S9TXxcrK024wI
s/NTviyeJsofO/wU9CCjmW8RnNPLUvZH54C0YjVYyngyblYRED6kx1sj5784Ay0lPJY4RbA4I0E6
IQ8CGRnyLDOqrGmEic0vHg6yBjSnouMjFOjCKhzfwvbkGY1W0GeZ0LCqQJef4EW3IKUV6IAYwLpq
CPt5JS5BezP9AhRlDXfrXTekctKRrnq93WBfWnxi8hBMJAMQod36+sOdQtHbd8rAwrdNpmOxFEvC
rrxr3MdZ/JyBZmV9hRV/LyBcpb8SgQI9I7Ddto0E7WUxhVynY4CuXh8tCRdqvo6pQJL+sZzyQciP
88hamHtRYqPxqMhRbBkgO2OPfCZsRZgOElPwNQJIrhxmfRxvJJIi3phmw7h0bmhA/F/JSYTtoq9s
MOCx9P/6qlatkJLMVGffnZNIymavIEGZzuJsfSNbJDTK4piRNTP+euSkAyWvu6URTO5tD+Icxeqy
UCpr2tshg9GbQyqXLzEHc/AQGVb45yPFpLHTxACUOY1/JGXcdPrzki1N/BvTvs/x6HDtvOQsQKJP
9XNT1/QWbeCLC/Jfe8E54EkjElQd/Zc1rgJwtQt8qyLFLp3EZ/GoCjSlewqI+V08vwl4Pnr00N86
1Kfc9QwlwNvmZn8izZO3bmijzxCkg2uvQG7sR6ZvOygFGgtMTmFb7Pfepb+rKIy/HWRptiwiks11
Hc/cTX7nKTykdEN2xpy/nsnNjTOT7QLqeOtpjo2JkjKp7drVOOadYoHE1Dp/UG+cRa7mKDlZhWJr
vQW3glmAxyzFEep7FIajjyLKU+qQltNtr3Lx3Zn2f22ertXkKnjNamC8uokqAj33fLTV+NZDyy4V
hjl4JIC4myJMVFh+oCvDe2miOzZVDQfzvVQJge/ELR0oc0iYwLh7UnNPIA8sN8I0FisjuUWw3fnl
DA5+THSVxQOVx82LTXR8hEk+u1UI9bpc/Bc157XcsD63bBr+drdJhVnzzzUmoMXgvTtRViKPJ5T9
RanQSvs7somh6hkbbYSPNWbBTfgwZ6xnu6IggiG7JWPKTdt7xMxIgmZb/XxpumKMtwr2UMxdzbxU
yCcBZLwH7OHQutBs4kx+ZTUvoU+UEs9fHuuXBUg8/pqrE+xO/j0GsS3d3FbGdb8JxL+x5LGkGMYM
iSJ3hBDlZhBfoMOiSClZtvfu+3IDV2qS13S+BgWnmK/3Iv0SnNYnyz2YiHcDDW5F7boW+gnkgaD2
h+sPbesHVEpJp2UENgQxwaokXPY6nlBPAvvrEaF/xU+daC5nCqmYTPi8w1G5acGQ3xsvUwMBpSd/
Hhh2u31MBYPySPpLBob4duK54188bevmbUtXpiHnBK9WnEw9H74ufCne3JsJhcye7CHNHoyBxAPd
ARO86Ff5PsOXv2Nl+QH5eMQ9cQVQuP+4F9Tbj4PRuGL0WlXDP0XgffvE8wDMcyMvWvAxIRMTX0+a
SVsCAhcDKpz9YL1EkNwCRxlHheenkwnTgaN7UCJRxCqyCOEFfp6+MjikqfStzvnzkhsaek3rEW7s
/VOYY+uSY5LsWGuszBUpztEBbcAJmuapkNVQvmVZCTUWEutYh4Dyup9/WdXQWNyvAttivddTXcG4
kCYP3AB7njigD5yL8a9r1AWULXRN5mfr4mA7XVRNaQw6rNt8pShaphQhVLfJg50W2fM9P4+F0Hp7
iu01ydV0XrVlLxEwm748qW/CtDRcSzRgB5jGg8l7p7Q7MRnqPm7JXFzfcyQJrYBA7cGxxgf1w9uW
MH6J1tE42TsD81g/dx8VWdLg5bqbuOJz6733Ve8BcHXMzZl8IsIHHrLznD79pMJ3w22myAVBc+cA
wpRUOgCrxC34c6xSMRjeOVFh8fysQKFYP9ULXeiLfdziz3H1jWZi8VCyOdKW5wAV06L3Ql7e1Mz6
pw7fGQBIJTVeK9b+diO2lAqBvxFHRfgv54U4pj7CO2nGIycbqb5kA+5teSqRrZtHeP87+GcCbVG7
s7TSjLkL4iJ7CuQQhtRXzxMcCmHhT7vZztjluci2FmI4eXitz5km89fUo1A6EC08xFt/CFYmdb6g
RhNoyMmQi21JZsXH66GBOoHwaBxVfRVgoJX6Nz/YbcZICJXjj5PneMHoT6c55JSvE4uLSoZmp+n3
pgbGDkGj7p3AVN9X+APBwOjdHzCIpXhT/oQgpvpEUdNiorIF7PG/9VDNJqg23WcLDivp3zQejLx6
ksSn8JxMe+CpWvzqVmWpfPQH1mELmU7V4mGKtXrHjm9ezWhVgN9dh6zJZO5Xc15h5FEibuxOjpnT
4YG6It+TrkE74qooc/OJGLB4qr+/kRofNWFwPo4QMp6Q8dHcg+QAEbdHs6kpCtT/Wjczy9z82jC6
FD7wSBqsPMgqmirAFesjUQbrOMUw9pDBNwkeMTcvTYBKwNmBMG4fAm6NLvsBDkn2peXVcxGd4J3b
i2L/x56rPMf+mrIb4oYq/B6jE7XVMVz2eeFf71Q8AYz0dHW0LBkY3lEuovALNrDzZpjvBVx5qyVj
CWL04qw2gyF3rHAg77b9Ad9WPWZxJHkK3scHDWF9ZVOZBIqdBCOKctQvIa4BOWTJN8o4eNT15zIn
Meubqvy4OvQicapI7D0pvTqt61YkcpJfgbrzOwqjeyN5nBs2Nsr63OUxmN7ZrGKx4CSH1YJCmxtO
4zQosezTtDvJy+4SSIbp2MwbwsUM4+8UsYr+NxLxzWKvjD1CKnW60q+F5/0C8peEbKISgY5R734Y
89lgI6B4Mv3mErORQ9tBfdo6CWBTrYM6oSiiIwtgnKuYrCED+6APio6ygGtYhtcIBUHa05/2UChv
XZe176GrOfz8ljKPaKKpD4Z5W85rrVIPsRorCW0c5Md3FSvv2a2UPPHcI8nC7aBEQvBt41akxCOs
IekQggjeBuisgmdSQCWtZIhwlZ8xMsssC1dN2ISEryuSHhZ0O0AaGN/vocqrxGyEaYsJH/DuXHFm
5sprabLGe3jY8Lr6Ssa1aZA4UfAhDVT0yBGHSX8LEcgzFEvvycDokD6im4n3/aiJLKLpxC6r8Tcw
EBHqYDMNwVC5bM4h5RlfBLbzPnj5ccHQmy18ne0gIKQbSs4bPk80hbgcfuDCidDxYOgg//XJUrfn
0PkemuxPJzJ9uKji4JPTASF/Gbgq4mzRKuFHmb5W8VIwcaHn0GK8Z01SGgPk4P/bNj8j5kJ5pw1o
Jx8i3TWoMoubm+KoJol2Hs/wBAyuhZccSST3lhg7V/1V16c+E34RRlpQim+2TxuMyFTQaAASwAbp
Bc/7bnxY3Z2vyE5wkLSPDagfopitceM2aDRCtNT6U80fuIQoxocGeolaPS73Gg3BBPWXhwBdIt7U
jWkX8Xf/CQJpbXEi5p2LKmcjC2woxZl0JlbyewFXfzfQjk9myXWkte2ts1m1sw9kgIUwU2JNAf5R
He25ucVzZmBmFzX84qWDS8i6NsOcJzKlqXfWR3Bgr9T38wpcye6LtkttJYcUpCCIhouTwce7gskm
u/bb0n/lS2VjhbodXDYIb1xTK11z0zHKhhPOSqNykcj6ZFuXOdKt1hLN7UGa2lkHsfSPNWMPw2cu
CUkUpyy9J/MK1Svy7x6vi/V3D07MatkekMOm35PtFysc3qkGwlsgHST9bFjO7YZbaxzogqQA8UUY
8PGpvebv6Bf+5Ow7PJtfq6+d4ruz1/+9Ohoh54hL3YQw8ogAOLcaSGY+2737lGCmisEA9wGDHOD/
NxFk0m8ZUQL0f4DYgDGQC3qzNmd8XseTR4tcMyuZZHb1ORif7ehHhPsAiNDwwatbeFyvYktms6Jz
kF8sbSki8rczZ/PaUIBVaZeHlW/K/HWMA1wyxfeIU8evEJuyqjK9A5dpH7MhuwDkuVEk1REWa2vr
LNxniQbJyM78AfsusTlP7yPDcZ5UngizOF9zKv43GIPUHU44zwZi3+UHa1kqzxxxPAPgh8WB5/xc
rnjEI/AwbZ4y4cmiB8GqxFE2jTdgBNE60uI/FJxt0ZMzNYUqSle1hntXn9aS70EP9S48SusHDQyN
E/5Q3EVQ58SEaewJTjXGJ5EZgzt7YJEh02LuAMQ3zqgqjLOA7jbJt8+OhJBrkjrIb3wsJmGTVNhP
TUBBDT/auYtHmuSZo6YXkQJq4bSK7+V4MkhDB7UdIXcf2qgQsntOtdFBXy5+ICFhm3OmXFY+y2Bd
+sppUgjAQLparAI4PZvLFiT1DhufQJky7q76nlncPT7+Vqb7jvZBY+51c4o5m/N06W+mDol8d53p
jlhdnTYU4poxeuoTez+7JS80MRDcgOVvaIfI08yLZssNh5128EI/1GYDXVKQ0KYb3HSQd5uWUjqh
0neygmrQHTpC5BhRD8wTQPuCBjCh5I/zOirqgn3ml2nEgJ2y73n7ygy3GxVJJzbYOzS3OZCHinSv
Pw1f6BpFb+Qh9Fm+eF8t+rocvSbXE2NPgcUq1AtyCxi23a1LFEfdBOuDgFje7RinG6YUwK9ZaDYI
ObtfsUVbgCP7/y+WwnvgW2/sNPWA6W96ocJ81p5HQxooqH9vaZ6IiZ54+fUEMhDd5hfYc+cDMWJd
AQN6axHz3zbb7ea4uaFLN4Ej5UTfEs9Rzi88IbRnEiM1OKLOB0/fNbW8ja/JYE1aCgTT4EDbn2MP
/K4Sr/VvFbtbZpZ6BhUTSzexoGGvG2Zx8A0dhv4UvZgK5tE0nsuGrSURXbPT3M1KLF0cSYjMnhlF
yIAXrpVDhLfj+VN9MMUG4JyFiwns8lMUS1WD3xEFIhTJp9Zo5BElScDJarIJ6P5mZXQWEiJrzqzX
v+Sb95zqWeWjnwbxl236CJn/dd37irEWavjYg/vkXdbuCsDXSoy3+b71PYftPBlUqBJZDNZqWGyK
chUR84WkU72wkz/vAtp9RWE5s2VkNUs6EvZJ9xvGFMGKR1wpUyPeiew9rzXjgD4cFbH0zD+ddaH1
bPH5U/zksYMuyWl46qrkRu+DumFlHanm+5b3sRvvZGSQSMzm0HD2dJBgEpuL/TdTqma5ORFUfdFW
+oCzqH+JgbosV5At+9DUVvTiCaf7ZZUbL1hbYS4h5EUVUuhDO7UU5NXx4MRaQ9sd6MpXMzINl95+
0KbMWl2Ei5RkbLIzMyBuWTp42BWZn5ZmTsWYP5HDDCq74IiED9qnWnNg+MGE40ZljHAtVBoELY8v
ZrjqNXOlmsXshcHUxWv8s6hadRk49OQNRFmzZhOcQrOpzPmiSi+X2f2hJoBTT+1PHuVeLw/JXAfY
+lrgbW/w+Rj+KcflbQFLhrs9ynFtetI9mxGA3+dB725teu7P6x/3ZnIxtCPKwAppIrfXKOcNuGJl
IVUobZhvvhbBcTQ+lqx7weRLj0k5A6iwUtzV+VscZ5lLN8DK/zNLr/hjl7yH4WQOzPPWuXwrMjTb
H9ULBU5cNLPnEEdhIGTtyntoMb3U8HEB/uZRW4ZLJaZYQ3yHOwBCLrPCvlV0XVL22tckHQ+HSHfi
y9KPj5b4QKZiv7Ru6BFY89bwL90CBLyNHa8OTqs/vb/eXGyoZt4KoyxjZYfELI1VN94SxvZzCbLY
n9rWr93JyarkuekJJzbZ99PayoR51D0bDZppnJ77jag+MtyAJHF7T+wHLl3pQyvG/G84cS0IYk2f
l2m5cq6oDDzSmRzMJp+2zo29mgNVoBobdcnu3+WtsZ6ij+O/7jEtyGRtC+UXKWYvXLL+P0DSn7hj
EMqwbjeaVeLjEmYGcd/RNg3GSHXnk5Lg0ghjkgzkSm12Sq7lNq5UdsLWMaTo/bDn6rl27GRUzPaU
0Jxt303/7dBF8qesVcZWdEvDd1jkeEKsC2TahTBk7jSvx1RXH3dRjYlxW4kayOJv75OTjflx7VVF
DYyiBPkgVibxFt5oIjerKCUB3Mny2KUbEsOitmCLUQwueO9IGONhMtmJfhujN5hC+/6FkK7vI4/m
rQ9Rt/UbyupR6pte7V5cfhdGThDNYPTi1mmyBFgezzVM6zdRmlHsLfZFqBipHK/qbq9b5JiGKGbs
j/rx1U3s2Y3+ggreF02cUGrhEDvCKEqTpGLbOBbYVBhYLn9+K9itJYYvnFo54yLrpDBtpYmpY7kA
NVIhkSSOBLAmonhwgTH05DjcTOo4xxwgn5SQ5a7HcASQoKYO+Accms83ngOKta+fQ1vme/vrln0O
uQ0GQ+BmCKqCy15iRVWxg0LDe/8MKdLHCpO3tmFKnRsU1EMzIUusRIzeeaI85h0Xc1+0cdBYtiVs
EW4yzEHO/jbVPLtaw11sLRE/rszRHdEzDl+nOrvr2aSzaMwEQkyZTFT2TQ2qbADiG1P28eTbwlEq
I1Tha4zSflbPgvgymvnITHO/zQcjbbNYZvuDHenULWgAKBk5ypOiq2pY/DJv3guOGEdwTUO+iHyH
BBy2AIY9V0Tr88sab2IOGa4uTsmHpPi9ZLcNt9QEUL92b2azhlOGQKFYBIqDni0qNHb0lAkKAqUk
ENjyuPxuB8jZlYdZ5LOI9fGvuYMmMBZONn4bMkce3tzROd9oU5xfB2OXpXooRpLUrAEmdcRbmf9j
ACAcX07b9G0CTsSaFQWuG43ss8O1sPZiMtW/OGK1OuBQkf17kDlgBzxUQ8Opt117eZykP3GHnrt6
uGU3KW90uH3XuVoyC2b9rEvwTQ2nvr1zynzjWQ13bLkHtv7k6vKPySrkMcRz0QKSXuAJFkI5a04e
zfY5OEQdcINUOs/XI945Vg0fiJxYlGOmW5yahLCjA7by4UWYvxePLCNwA8GdJ8raeoaxysPBWMvS
tlGfCrqypk8lPzppQJYIMVtag6GB6iLFev6ZDPRKZq6M11irRu2/6XVMy9LkPSdQKzVdhpCsBuHO
Bxi1Olctjf+TfhQB6teAHccZx+iaLiedLHXBwDXD6+pmsLnnD+eztbUZ17YJencUHWUNU4zRMnV9
BwkoxdBiHGomHR6VoGu7BHQKzuMaEL/9hpk21eNqwEOMQUWXaJ0RIDGCecatcyTkWgI5QtJeXEBI
vXB9Zru9Sb5FRavBmia4Chvj/+M0LenFC1WcapOKQ0Hewguj/gZm6T0UPD9cw5stXHNlq29tgsRb
/cnIk3gwR1Q2++r12JYH0uXu2OXUg/Tl66kU2fPNdQ2NLyQNE80NTSpHcNIAqJLMyIXbKha7yoPj
HxpQzR2gxuf7vtbl60yMIj9f5hhR5gD98QmbkGu124Jd7xypYJYvL2tnrRhOtsBESgGi6OzYJ4Tg
1KeVkF+O3JS3k4HcBcVj2wL6XxfOES2GK6Ff86PPoodhytaPvV4UaIjCJjGMK+XNZEYmSdhPGKiP
OIyxVHW/o7ZJHkSnesBvsi2L2HirDooqAgFne+A9IuqrIgRJ31rYJxliTH8R9pTxpSAYFVV6ENju
7L5NOJO/MWjIemhP8GkF99/xLVhjmXR64h7fzCL0iZJH4E++/aCyZVjaPe0ZXthZdqpc1vapJC+0
8yVMOzpXWQ5SPpt1i7yrsiyzC/4Z2yXgkTZPNjNTau3oByolQQSu2sRTBHYcq44tjQo6yIrX/j5+
LerHKRbnZfjaLketiL5r6gDcUFasNm6m1xOFWCobXlhT9+0O764h7/xs1gWXXlvZ0gmNNq94MUss
/ct6gngyODtrCf09faPPUOCDBbjktv+kyUSf979eb8SLTGnHldkIzyiNY2mIAkke4OWTS3PfU41Y
NrNMX142LHhnP6oPb2vgQ+mVtr71qp4Cq8uy3hGLneoXuGoAkdNkr/BEwkWmwiKYatoE6wlB/uGx
SX5XIHJqMoz0rIodBw7zxhraNeCyVBV1v/k0DnvjVIcFtdhlw7Yj2079WAqM4fibQ7sRRpkbgq5I
n+y2WRYf6BnB+PoVcGyVe2a5NHLBJja1pITjh2hMwJygTYnic5u87DXfT5aNi5rzJ0INahyaCf1B
aG1JRN5jdD6DZxDVL7SfEuGij2uBuDg0ogP7aQJN99wCn0/oXB7vR7k7Uev3Vi+TA/4QvC2im6Q2
CeJpotcMPzqdu/YM8h4iOnYu+h67JEm1QdxLBqhb5GJIoHSfbcs7w7kQ8EGowpGhL/3/aPK5BD/4
cC82CIcgbdr/811I897EUuohnynreaaJg+k+SzB2ZZM7YnVNx0Kq9k0AAeFjw/ngLgde2tjRIxfK
DNfR5w9zpfOlRS/wqU2yozRnhyXIn9Z7UTcsnEj4EvMfR9W3lfcF4yWpIj36RivH7qPDlPhzoUFf
0y8BHsuqMFCUX4b/8n5no9H2uFFUBLoJz7QpaBv9vy1qiGpy288aMBS7psm8voJ617yYdzXLr36Q
gsfCdUBbWM8ztNDkz980BZgEvPX4Rp1CblAMGJOiK+RTcCB+2ij9muoGz1YhnO+KrNah6tALlASx
q4UARFBfhYsJy0ItZceVf+ZLt89FAFSters8nbJVWfR7UFP1UERkZh+MARmI8pLOsEZwzHBpHGg+
WMVKyogCVdClZw+SMAHlr+YHLvgz7hyVVQrn/lrAA2gWr1nWzcMn2aA+tRi/U7Q07b4WGVOu3y/j
HjWLf08ydK0Krdm2ip9f+BPqo8qrJk+QQ274Cy+5goswzzizGfpBV4vq9CfuMfesFzZNas0Zo12t
pMAswSJOKW4RMU3Xk2eWVaJ9douUtU1JEb6+E/IACGSRBK7Qey5/oqbOMb35Py/OdVTZvjfZci1U
W4UxI21WjT2YMITNOtNaUlW+tGZV5h1PWWSO0mKNDfvN5VOJ+Eb5wvNCZnAm1Q9plrb+qM9EDFHt
C431xcWp6eGI+rDX4PFBMstZ1qeJt5++yK9cK96uZhp2KWdkbz2g7ssJ15PDRv0L1V9rF7F9XAg9
i4qVBR28wL/OjHvrDjlbRgCywm50Mg0UDgWanRdgK05GYoFNoeRc/W8d4pftRR6k09uRvLlWVmqt
rWuBCJZZNANIQaPFjOLXzHO7oe6THwwpapbDmekGu/mthRkrpLsZN0apPns5tHh23NnXdoixBo5D
vd2ajKgdLTTHVK6UtLa/6QcdVRlusEc7qjyMMZw6qhTp1/r3J4C+SSl4e1dLp1PdSVaLJ6JQb+vM
uzLLiFZ64/JKQUd5AaNUOZ4d7TeGnu9E9Bfc9ZhQ3ifYM+VeMFhELnRLt+jIeG7/3iLu7PKHYdXd
LJP7fFz41FY3tKAwQKQuKwDozYfipLW4Y6jzXXTABGgQ2JqJYx/MjpVjlOsFENMsD98VzSsRAttW
74VKGHm4KZk6TE+VHjCHPxmFu6AC6mh/9v5zdJOLCgAJ2g+efRUAevNQ6KrqR83nmGOiBlMWVA8s
8f8LhG+RIbMjTi8DrhTOkvctLG1+yGpoXDhCJOwzbpiuXcRxg4h5dNAQYN17LGLT8S6WnyJSD69A
mwglBKKhg1Dh6tG6IneScQ+9qf6zbCBnpM4UL1lZKL5x/7W0gxP7zPf8EHFjw25+zQBe94amKCRK
vAQgeFov+KMdTm6SSnrfnKh2ULVy03JIVqR3Go3nbyjFxiUdR4CF5lcH93dG4QkLBZp1yX3wzaRd
VFdd0xseakWy4mI2nygb4e+b5oJUv63naANgtScx1mDQaQhSLxO9bA9lwOiUKZMtbmWGnWqVX2/t
iyHg4MremPt16GB7Kqx8jWWTa6+SiV6BSWznihxBpzbtYNaA9A+EHAtf9SNK6Nf0I0BK/04ZlEey
z8GRIpVs52kY0vnPa2WgYVoGWJql7GT7CwPOhDVLWnJsoZ2Ta6+dUzcEgMz0jwalYELqn96EU7sJ
KUZ/xMX1m1VIkqSs2DvdE4rVKjl5x5D/p9GjK9Ub8M2mzNBx+Vm/rcIyb5uzoTGFLMJqnd9AO4UN
T45J+1SyC3QFdAikFdhxPPJ9NnAR91cIon2sChxW7xka19rOPPlHLAxs1DyNa8XCYc1BQTb8M/7p
GYnladvS72rJJiUyRLMDb8MusKPaoH3U+RRbqnWEWXoxgRRod2ytfJSSG+7R7cXyqIBddrioeVpo
0BX/ZEMaH4bhO/K4GLR2G+sznNE+h2fWuIc59w5gRQlcILHcLw3u4T8P/VT4iiGtNl33z0vq9KwB
wBLosnW6DjHrhgrSY8hh6L5VshmTLOT0k8dZWDzVmNkUIPHl7qmJUT1H+xzlvKoHm5uE6tvSkcE6
E9rsFUugdMsFqDWIjR845YVLdR3004Prh9dVb7xwPwCEhRjT2rK7KEYU9VdojKt1j+0oLbXLMYHX
QUzrRoq6knyXjC4G078ROG1iFXvDFLvPZuhNfDAIGWD41Wc4ZhhcG1uXbFrpwbK95kuBw7XFQptb
tZ0DqJ8VwxEqe1op9MDLEARZQAzfgzqL+nGro7uTcsHHsmUMY5X7l6a/CDQy51TV1aQnJTzfyEQu
rXPFcGQbCVgCIjkrP7R9B9mvvb1la6e1tWOqeaA+LN2s8w74aKiaQLC6BetlbGFeZ3dh3kzXo4P9
gVw0XKU9m6FfPdmULGHXelFiiMLjo7UsIEWjuMAnOQuu8wkJA5U7vM09GzSKy9Sun+LLjXwOUT2E
jSgODWTlFJkLltp8hYCYFFGcEPlYf48CLx5eN2AxHViNPQJ8vcF8Fr/bkZ8agXuTh03zQsQEJfgm
ELI6kfbCMSZt/km6VrPC17Q3cwVNs4vQuchBgDuyNl7r8n897RMvF6uD4zS6zmvW4zHIDz7JEAYk
aQhSL6Zy7deWuTN8OazzAyv0Jps9ZaEeX5dKH8psuVkoGiHqzXlHWdTLeh7UD0415M7CsktdvnDi
q9ltDLLAIVAJ83nhFE5UWdX54f0clqwCbpeq0D2K248Z9zJ4suec4176LD4N08tC1tpsboup21qZ
4jJkw87DLt3syLtZJsSSRzTbwN+996BaNAZjPnDOZKtG3q1V6fzP773R8S95ytRLfgWmqoyjLRo0
u5X8b1Im8LWvACFOZBQzQ9jRHyqViiy7BlLW9OuABf0mN25kfATUc2F3EE/8xd8jZDnD/7AVhOga
yIzPnZINTHoyHPW+FtlKrFMRsxWI5QwR4xRfDrCsUr5sP0KOHLr+Ck1v4cjWfk4V8lXnBwKd5LVu
sDZzrjQgrz07PyqKgsB/p5HfeWE5MDfrYO9KBD4iKyRwPWzaplxBNr6mnPp3LzVGXD2rjKwBHm1r
uJZXSgA0PmyYau+OOplFrmG9XGz0HreJJg5Zxf+nK51HnjuY6xamQSmwcvtHn3ghySoJ8FYfFQYu
G3Ntr/elc8h7Xj6S5vQngIcRBevanRJ2u6cKIV/RcBTp6ibRDuu1ZpugcuS5h7z6IM3TGcivLxNH
JJfNGbjFv58/wCGX+ifcpVK1o38uVSOpLs6AF6BSjpvVGu6CgleXb1WZXOhNQwlyBDEIgy/9thXJ
BJ2q/iRtd12cneACiFIpE3NQaspa9Qhur09xwu8gHlgSo9iGLLemIubSpzQ6+RzIi8SQNhx6nc+4
yxI5bkQAeKOidGk9ZPRTW9GKKxgPRqpHJp6s0ZcOLB78oIPFbMOZELPs+U/Ph2TJ3aiCFkbFM/yP
yFpfgezPaU5czki9b6pnzOHkoogwHmM4n4/ZhvrIaFc8chLc04ZzCbnESIA9RWHw6MeCipu5oCho
AhlTFJ6pFDOfJ1AkR+8P8KuwdpkYiMBZltGQxRVGmuDyS+yExz/taWAwTtNdNmLBtGBX3rsgvQ+9
mwhB+5lgvTEcgMzJ1yl7mQJgQ8moQJsz/KN6JJDKtHizJMaWxOlr5krcDq7W2nOQsknO3+qovFxk
c3m0P93Kv1ePymUNEhB1HNeSrvLgssa50rYY0pTB580wW25kD04nkQydOU94p5z0NFyKicM6wc+f
tQ2tIUh4ld6karUMhc6jTDTJSUjN5Dcx2s+q3HA6f/sfdBhS5dRNWxJW+yGPtYx+NvYPhRixC+5J
9k4loSufuKFkOfoegphy60C0SC1COG3qYHreqmClv0KVRAkFVUsK9PGPIUd2fydRtBDtRD8SEOqN
EDSSOuTZoDdtCUlKdKBAuk+bxTtxTjxrIaaG5S0auI6OT+U363iPEoLdUeU8/faFuTMoiNe09Wj1
Yp7zblThryU+AB4ElkJ6xcmjxe8t6E4btInHVbuviSMUhfLOk+EbS0ND4GGQZ5Q4oh0pV3Hs2R+0
rkWawiRCulmJxXK2JCB1h8fkOm6SaEAhVXQVxhdZ91FHqlDuyUQRIbl+I3sJqZGwcDpINAtB4ZhF
TYj5+cXwDmROF0msUKvWtC9l3yecclaOZmmSIv+Jnh+O412CNfeeK+ubDtLy8i/nZ1lvA/I6Zsg0
RWPV68adOhcb++KoPG/Fx3d8fiSr2FQfcolGa8AWKp0QUgwBSgIvvYN3A6Bi5ZFf1pKYBch8M2/8
T1f9UgK+B01UlJvNx9aTI9ZeXEG/VG03C50XCgAsqPwZBKIClD83iVHi9sN0jfA63u8iSSYQVIgI
TxgauxtRSAGXa1VuOJ1jIK+t9A84ijQljKEx4xoJDyhVq9h+W3klD9oTSXBsGiPJ/DZGfiif3mk0
/WirMGvwXaslgOc86HVNCGko971c5RaJ9l87l8G7pt7apCYvxCACwdQ9Mwq+RHTkov5nWXUTALAJ
9OYmLR9r9+671H8+1UBujmNTJ7mqHQsx59rPW8vgR7tX7T+28blmMxzWittz73FT6SGRDja50pJu
QltQVq5C5QaXXpF/KzjhyChpoEGGp38vUsQUDhuAycZlQOe1UkqfW+s/iLWmQBN0dRJxLnXksr1j
osg8hR4Eyl0WBptQJC+7G9EUSnbqb1ftTrwSfxx3Jt7tFNPZtAaXdJCbC/c8au3eEMq9/2hK1kxs
pV0r22/ovBxx2zvIWE3g1LOmus00hlwYNT7WSzj4f9FHMjvJWeZ0Gehay4ftxMgAVAbgMQTPXlvx
Xgb4lgq0V5Ihff2XeRNdD9vfb5jzXXFqEDzgNhmP4yaueN6+B/wHbIEOeoeqvrq/pz23Lye5HcQO
lqPNBlsvfNz3UWuzNR6kHomOPaoE+rthFkEamn4j3nj+EjtogMI/TlrFLHXxsw8PPwkmJKG6wHac
8GAebr6lBtvDT7QcMnbeINT0jFVlW6XjFltbUrO1Ml3iTEaorWSrYWtxN/yrEvFRX+s4vLqnN1Kb
wKojEgUlLZQIaO2hudSzC1ZLF3kJ8gY3un14Yo37A041uzVmD0CkdaxYLrqeKbXJhuNqTLsX4FWN
XuYBMMmeCmgrOZ6JB3x7vxniI4ZsUOzxN4ooiWcM+jLflT6Yi1twcK8868tllFlt2RpdPsDOfg1t
6SDewYSpPdXVB68knkh0JE81LNZBIPcoaopE29vAoPS4pImj+w+j6QGoHnVFOxkb3uVsjsBPHOG6
KCWzZ9JKgOvgU8lBBd0+Z0XxaMTwZtWP078OHhPnu2vjjcE6FgdwU2/WVuORmLGITufazBZLBqyO
cLBBv3JqW1xP5o6g3Dprd2Hc4KxvB7QzX0psn/L3AFGEuPWTZza8+c8RwDZBXYD/2GwK6ltSsuNP
taKG9vIKNhOd+ypssm6N7g/feHRUKLrWsH9D1c9F2oZKg/9vTYoazfWm6TR58bm2V/ZBLUx+pHUV
V6hcl8859fkKklldl+X4Ry3DRcoJepGU1ACmUOXPvO8B9AhpTTFJV7CdsxJmkWP/B+kep9HQv16n
5Dd7CEC6woD45Jx1E1T9xnEl+maYAQgEP4edBEKnP/spe6amZW0nkwb8wQKbRC3hmHc84jE9ze5m
p9rE10Klt2a8zlmDj8GhkT+jfNpdd2IZngnWkGx1lxKVd7n0DIBgnetRvjX/xJZ0E/oHGduMHd/G
rTan+cWxHtEDT88dI/KI/+ZPAtL7j+wt2RiHPyvwjcgdEWkiP2ZN6ZeBD5weo5X9WooXcg5M8NjL
Nw8yPeNDODEGyccFDPOhpBcu7sxxJLPbvbgg+ZzpcI/YnpA1wHjCofyuYMlX1RhP7piLe5IDVvKL
8s1JI1Oy/lcFNpE2o+ZAp28QAiRkKTuF+RGROd6GfM9FKYzOSnn0I5aPGeQsLLznuBDGMVxo/OcN
x2x4/rl8ImvHbPgGj8kc2l+lH8nRlirpZSL6BxkJGKybIzAQcSvytyl5/joItHOoh9NWczss6N0W
YYVdVg4stZypO/Zy4/nYMmVw5tnQgOkWM3dwGxSfLpTFYp4RcD8wHsOgdKLXeovslC6IfPSUtgIL
5oHKOUayurqr44SDVzVGE5ta/DqYbB0NvFwzDVM9I1JgcnS6eSHdENwftrQvsXqwBHmZVa+DT4dT
mlPVw56Cp08+H9+ZP/qb8kTuyp4LYlbAMbyLF5TUEHBDc9ALW0u3QNJOjylXH9HiO17ef2bliSeP
vNv7Fms86azlg/1SuYHbO3CdW2RGWIhT6eEz5d1QVs4CWTO8X7ff/hE+FxWGGh3rbOOYp1e7F4C2
pJszthscAE1cabSOHEShq2K300yFXehEAxtnM6/ga7WF15KOUsoVqXykHI16fki/LpoFslDX04PA
291aStKEPA2NikNFcnRgv3wE5BVy/Bm813jzQ897/QKeJPcYFMR1lEmSGukQzy99vLLPvrEsxijB
sAzdunhyMb1y8SQWM3ITrhm6t7wcV3+62ywH05gm+ma56HO7uuDfKqgNkgUMumQClZgyRWi2a+wI
9YFFQ4adfE+aKvQakMosQXMpW3B5LmTaKKNF20d3uIWHwhbTwkoYjVHJ7qXRzhlnywYrYP7E76JZ
QUxp4/9+pInO12m6N6QHkAKVWdvAtwIgqdOpcENQcQ9kfIXzluxORvarJNzcJ8os6fkS+gm9hEXS
qNqtLqKWOVYzFnjS1QDdFp0MVSknBZPpzhLznhqjGMRhuviQ+gUYfT+5VT3uCTHmy8v7wV//vD/Q
dtXdUMXiE7/9P/IVXMsCWKKoguf/zsat0SNE+oO4/JdAv+3mOl3Br1tB936Qle2lFZbxvY01didz
FGYXwHUc8w4+LfbcPDCs7D2AyXrHctXU9UP27jxz+cHFT3QPo9o1n7RzHYBuQ3ocid3iDA3SdnYQ
NvCubskxCUhE4xnU0UuiLHRVx7Ic8vZRTAE2TIP01GccxvrLFz3uRhIavSOo0wy5bbwW+aZZ6Ix5
tVYhKGH2x9WzaCdpEYO+FfboHo7NtDdFjpmKX7g+4NxQV94uG+Metw9lxnqIwO8LYbH/SB8SnFIq
PdrL34ACAYARuOZuUZ8JladdiUDoGK6N/DmWrrFx+OFU6YcKUXnfWdwPjPZtYQGVDyeMjYPFMXYG
Q+lE7zCBtaVjREXdztIhYVtEaw8sn9tNeDefPnDY1g89ET08IH/pFwEMGStJINi40ZcSPqlyXPME
MH61L9dPotcjwVdD3kibfQiDa7BPpFaGEmyqg/Ty3a+f9SLL0SZtetpa4FH0nco8K+Jxfie0fw69
P9+I2RgZEilykxkxyXVVk/OZguYrHGp60dF6LteGpocKRcx9JrPUbkDKRnfOx4xxVVxKeDvdeQrP
MXdfJ6tWOl0X0ukbgOdISp7rXr57oCNGnuZDpIo4PjEADudhcHuCv84FZlsS8atGdW6iLVsBokxp
0gQMRLaou3RGYMFQs8wKLuDlP6lmJejYz01ReBEBpWet90wiLqsQucCn1pQloRBGoUDZO4vsX1kz
KGyPzpCAs6KJpUVfMyvM5gTUhKMjrMU+91wk59zPBC+mIA3IPDy4aUgUfwnXFRQTHkyzPK3Uzd0t
fbH12TfAFZtluvBDoZMCQmTSSYJfsPljn8MRBMB8yDJIK4fZXsxRNP+aCpyhsIEnqSAQ+G6OUWt/
z72hn8Doy6oVuLVyJBUY7YW2rttMmqMw/LnmkVrQ1maCfQ8ZlruJb84SnPZtGD1ZDUZ88sQSRBib
nVgk+/K5VteN6brA3evymvOFSfO2KvRu/RWzqfpSXx13ZQwqKBOjxzr2DhNZSLPHVY2tPRfIsxQN
2oyNx2wBzYBsRiq54t1o3K+nRVwJHb4vKsleh75q+ZavlMeNZhGqS9mMHUj06iVOpuXpqQj+BUg3
CS4qm+m/cRN4IVF+lXOkgbV7RFfZq8GssOCgRRQrZp4QDmmXE6T7UWaDs0bj6nhr9K/kZEitST3x
6qsMBJMTzo/kDwoLKbgGbzA5OYQ24F6fJbrEidqdZisdwkN5/OJLxNu0MQiF53hJ1grz5jVlWe5z
Ig+anJjL51AlJEhqe0d+B9fit0Dw0ZLpREK/mGF8c4OcQ9GDIaaB/+MAjPDWs/ljbRl0Sm6M47q+
5/r/goZo1QdhJ5oGfM7pOyXI2FQKdXm8U9s99hO5TVmnTd/sDIhppJYACWL5jjLy8LE0hJE5SBWQ
m+6+OPcgHF6EL6Gqk9Q6zrQoVXjhCDmlssPl+lru0FVspF5ERaD12ykU3uzNRENw4tUcIj5GnNKH
S5EWa9pOooHsDBoI0vtD5P8j8FrswYkoPNK2/QaexRkna5NZKoxKI85ehktmSLSNVQBqEnJHCM9f
pED6c6b8OLlUOjZOhV9UAcJZcG+LrXQN8mggKEqeyP3wbonQYb16NrF4BWk+2k1qrj4RkNAU5Fs5
8TH4Ja8FbXBXw031aTOaSkOwZcUimB99X8eh3d7NNsUzN5IVh0hBvyAzm9PBcZhiI3R7uc7nw8DB
JXsNc8JDyewuh32zHz5ZQ5gCCH72e0ldAWBr4nySJt+GM5IFAlW1q4ke7D4FBQctUSFBaf+AAM31
r60bamZHazagsZYvTZ9daiKDPFg4ungl0vFWi6nnwH6zwLqKFBGEAp4jpqME6f80sN0lC2fF3xlg
W9O7tsJfa75ypnKfYDrUBtuzLTq6eIeyZGucsazWTISLLK5RpnRw86QDMLDoidq1qJnknWM9BdbK
3Cbvs33CQh+VH9kswJ+NsrtEJAOPo3eLiuuRMaRt7yJJdZ/Zk6SdZ9p0EXkEzlT/TuFyn5F8oAg0
mjASselNA22SVAF4pKG1XO8OPrLHr7V/lAV7/0xF0RQVSgMOF9GcYw5xxaHi1odzt7sl3pyvOId1
Px7wje7/2PCzG6eD30TS86O97dmOey0VsOdjxUwHwnR1nYN7ZnOZ2UhBlGDNmPUwEP7u9F7JG60G
yM3+JSgwirsxlPPyNrzKU6Iey4SsixTr8oAFHN+3guSgWyXLoN6qOHHcrW2w+SYqVWdmN1uTl2My
lw684O9xWjEZrxItsQakfRCbRwN2DSscWFJt6alohMg7XVv1A+Fwv/WhD2Fs11sBJYaaVSmjp/uN
51q03jHlRnwfmjtDb4Qv1EM2gGEfL44aIOuvg9QlaV33iw+XzuzesNYOPdBYHzntHDXqYmVPqqUy
B+jCfqJ3StYzmxGUJXARZ2akOwEJPAmVtuU5jGiCDn9aslDwT9ljghoNhKay2/HnZDUrdOyIyx9u
zhrQe1yRJBhp/d/6yx9yKN4eezD3Ofg7T35YoVtxnXf1Akh4398uIoae9Z1sRtAvXtf70m+AH1W0
swcleqJemSsVEMQUQxUYwPL+Z/59xdmOX+v04hvMv5BAe+mz41914/yDyU5y1TPgIUQQI9gL8Jdi
PAVbRTopF3RHJmuWjtgToWvEaopQg9+3LxymYcrFIoPBAlb25ODYq8BiEywZSY323D+TOT24AjQL
wBs4XqVyxuRSSGYfFrv+6oLZ7EHEUnKQkbezZ6E1jgbpax+U6JgG+358SaeAgx4B1MhRmxqWvqb2
F2WCSJQWZ0Ug+M5srAemRGZz4D1jngdujL2nmonXRru4j2thoB9p0nLVvSfusarWkdi/yHA7TPs2
r4PgOF5LcWymjzzNm3x5GLdJ3OFiJ7CKtQIfVjPxUdZvkc78recp+7JlxoxP7pV+uYmmVWuTWO40
ZzaZ9TNTzVy3MpOh7TylxeWNw2Bon9vTtQ0QrjyKabiPae8jN7V2zclw8R3kSm/xy5PYdUUyhPa+
V/hGVZ6xtkmj6/KPZdeQ+xZiPFtTxRV+8d7oNEG8yC17cb3mJgrjzxPmSz5VvyNGnnNi4YS2cddi
7421jypliVv5eKkTaB4ol5hUFAsjZjMAhTbOlNRYXBhr5s+jHN2xBdwwxyjZ/eKzoWJmhFwCfrVU
rLqlwZUd4hF2E2ZfXv0Zkjlz6dgYtmsLgvKcRG7diRzG3JU1JjXKSGPpNYGwiP9/xMykkK2zu2DX
fs5EVh/A7DcT/eYoXvpjuQHG7GdbpJr60bAARwS3WlZW0biFOoXM6AtHNJgZkQIS/hFsIB8vYMBd
gF0MgcjSEdlTNJyzOP2hs9yKhVv3UV7RwXj7tg9J961eQFnceJR8Af68megjabeQWifpMme8g2Sm
AEQmeH0m0CPpRSUYSkrRIL+Dy6/o9gJDv7a6B4Xp4dqWjN3dz4zF4wTsngZM63TYGY8NRK2UPD9r
BdUFKcB0ioLO8E7eKeerRtxEJKH1Pa6GhxHk0GUN+5t9J5tDpxU2xIzTWONaLyYnTge6zF6mRtee
rqIH8wIVpwVfcrCj5WVwH4ntsIPi2eVGMcxM1gGtVIZr+luMLFNObXeLqj9fq6twaqBqx5GpEqUf
0s8+zGhx4AcqZekBEUEQFTbFnNW10wkSNGds7FSz+ydDFuYIX4TQ2lC6WWvOFwmLedYUkKwhAxti
I70HggqJJuj6tmiwCR/GN22U0K9oUG/pgTyuPJlmdf1kxYPtPF38pHZZehEN4JRalReOM57gJe6o
1JGJPX3IUCZK88YaTsmtrCfyhi9QNS+AdVhAjcVezAzqBpPnMs28i38s0a1LKhc/bVbfwelm+nY7
TpdxE1YfTetAQb2ThA2UpDN8MGDZ4yyUMswMbRhOcTNsjC8Rklpn9M08RxQmpZ9UZ6w593jfpe+M
IEiERofxfyLencOQ4XLWBznzHspHDTlgaFFH5sj7SEaWgUI+7cs9yIlp1n2PpyW+9692U0oEHc+H
MNjuwHE9eQASdpiBOrhFePIqB/5dQu4vVUsuakIdiEOA1HFmxsaIxNwKSqMWAiqNvQ0Gub3PTiU4
AepeMVlJb6c1FCiB8G/zoXQUksrJjKot5Ypp8zoyf5qtZyqttSaXUydIfNdKbBSYMoWtDG/WAPXU
Aa5GZl4OG75pjOKXGjNpAqwzoNoapq/Lc7jgpHlKkHAP91ZU+ibmjVHXyzfdxsHekjaK70pLSBdX
+kEng5zeBUVOrFIdzno85iOKuA6WapG7mnYbph1BhtuLz5e5J76nAWmlfJ77axPSNPW042o3Yc4h
og6uj9ZvHmF4O+K7n0V4twiVkarr/uoiokWG/p1YjyCT0CRdfYMRl9hLhyx6c+cxjErqoTtJLJZa
raQClD2iMeNaC0zWvpp3U7J9a36RtP3lkFMrfQF9GzwYd1yOFL3e9of0k9Qxpesv7BymtafIopgG
4VZ2Pdkic46K+2ctmYyp/9z3qZWIGjEcn/uD9McpGWNmBE7r5dSLmJIz5W+rh3JMAtbOITLQpoXQ
oDccah8+94T66b3ikmHG2ngJAwmqv9U/O7QURlIJETClPxpuNVjgxQfZ8wKOzLmsSIIEqFiWG/Q8
M/tbiazKxWWgMpxay9fh/Dq75BPu3+1A8/KfplYqhcfVMak2ZALnq9PXZ7/Brh/DaDmhYZuMxafQ
NSoyC5T/T7hAcI0vTZx6JizQ5ZzEbzLo18eietD/nZpSUO13li8W9pNwhy0Rd9nSgbbMT+3PC3LS
bSavpfvRux2PAOMtkQbE/ty90NkVxri8t0Z823WJTtl+aqAhv3nHo2XUprFgeyWOHHBcNvsNYrKB
MGKx+OLgiAk7hNSoYdQoNxrNO21tXe1Q4y3DN8uADI/HgO78pNnobT1saHzF8kJ097fI18Ob4BrV
1j6HOY9pNlP2dOYuKe57ixxXecKCWD82ujKcgYQWhECIsJaryiAJEqruWkAVKsc2EvRvzj7AXAl9
Ikxs9Tfp/iLvagm6yiTAnM4UBBlkJEZ8KbR0XtNCiPcB3qn+0g+u5sM6WNLc8bK+xDxM+HzgFk9U
RrpHt7D/ER1b+f7yqzmg2vFNIfR3RgfkFrdcyBfp2wTw1hsbkKGv6IPvHUtk2ktwDHKVbCv4VWwe
kTvNHHBNDiTLUgfadrjwLuT5Eg672DHFykC6C0N8+5iX2yc6SUpWHcYQjqILfwhBq45yKEWTsQOa
6FpIgkKC4mp3yUGoyK8GprwakacC8th8GnjHevCDVX+y01Y9N6S2iUsI7iKwm68Tm5g525ar0EFA
GlTBaJ69vfBycP1GzcifGEu/xib/LmD0Uaaa6XT0tYv2FDLbaB3hR8grQ86c33pSyy8cf1HeIcEc
Snn/uYbUUGeflucYEMtZ9FS4aulLfWbdzkXj94HmIItvVZHrduBn2Uvt4fLWSks8ufL5ksDFNyuh
yQLgCZlUUUjCcn6QeiMdk6jcxli/phsN48E/1SjWx+3mHjUjICyLCsbNCSaeXzQtKobSqxIgfxrI
9DKSPVKD1jTuXNJxAqArkdpUxdVXIzTva5+yLo/yTroA3s3MHfORb6vyFYwo9xCpJbsMNKE2dAlB
tTzudqdKvXZ1jQAvyz6UcJKZ8y13ly6UYpeF47Fiam4Dc+C6vheM7PSRY6p6FCmmZ2DM/IhwGbsu
PdiGGiVt+n7YfQBCZ3rzkKVpzy6QrqPs+CDpmS5Bzw9f/dy23yjOZJLTSGMhEQOQmsxhWhUMNAiD
gWDvLUUipEi9Ns5Gk86svEAP7BFaU+ePjb3sWwoAaUGktp2rWQCFC7QLrlZ3Zra53mBpv7UwKlju
P0GVzsvigvKummSVDmi3lt6JsrFdfOgtPpllygpX+3pennHnWH4gf3l1Tn5HfjsZeluXMvN6x36n
3RGtI9lVdcrZRgUYGbO1YqWImTk0MJfY4v2gDNhxXgQbzeUHWo812j4pPJ5sQ+1AtvvSRzPjfXbx
pvQp9NPX4nHqF7LIYfMjtiJ5MPNQy2v72rG7Kqr0ueDJxq+KNhlvxNlruO056oV3IVyogD7A7CHp
WJn/lpp81d5pBDkc5MxmV6QiDm7LOPSWIpd+w4HgAfWrS+q0Iagz+noCFa3nz+akjaIK9EMmdxxY
ny+9iueUWRdt0Nawkgw0IpnMdCAq4hUrZzq2761jzTm90u/4E27BXQu+oN5X4Jb/ETd+XnFX8GKD
zClrKRqraUopslwbalpx1JcBAKidLF+qtDq0IaHiuya6Qb/kPFtgIDDsj1kM/4p8sgzp50i0lJ7E
7FZU4FJdSDl3edmqduMp1pEZIPskTKHzvMg5Moru8A1EQ/z9w0QopwqBMji1xPkXO9rUzeGAA24a
9bkQnS1G067Pqv0TF4b+pf4PgOlySrvofONhZnp8NxW5zPNiXtNalp35psRGAxypg34C7Xfc8oNl
ljBRKdhlusWGN2g6oFFAqYQ+X1E67y59PEwFEUgzmRJho8p8UxlBaz3Rt+s2VBVgE+vf+wJnoIjL
F0hNl/ztbhjnf/RIKOBWeNMtpfK4evUA+UOpV9wgL6L1faVBTizL0iO+lCaToWAtOr7lQc55dy3R
w4uaM+cwr9trsTQSw1lAYLP1D8pFuxgZiB+dskiETSH5NUrAl1k2GW/Yg3pwmRkyvV0vAHB8vQP2
rmhxvas641xB7Nm1OdqvyxzhDgO6lDputg7aFMch9OW2FkLgW9Om/2PXh46DaOEoSA6xEt/nh1Jb
uHNOvjoUqfD3/ulQ4evnxX4Bc58Lfjg9wC/fXXLiQXryATnmeopprGX4eKTnUKWWPaSqh943tJCx
P3xTN7pjExLkG1BUZ0DsrOS3aSJs+0h568jCG5PuAf4kIrofVclRxSSN+8gGwS+d9C+79P4P0gkK
SMHe8AI1aO9NptCenQ3A2S2Fs4iiBoeGSKqTLpUX4TXr5l3SnKS23A5N7luN2jrZSBNVUZ+JAwTY
wWS/9xoJmNOZ82cTZwXWpeZa2awyA+WR6i381Q0wQvyLnMPMbPLeYpgHN3c5s00dIJ6e7izwn4XQ
w8rpYSRcKl2qlvsEslf7eryLp9zxMlsbOgKAKFNDufhoV+3m2IW8N2LyHegl86V08Jm8sOtNUwPB
Dl9aGWVheKChriEKU13Sr/D336NUCmroAl3i6njrfMgBGplK4LnUb1mFGBEA2zf9m5ZNvOsCSiR/
5tO3QDLfdlDw2dX4Wf5FOyDTe3D/bWocerz8NKtqQvvTHnaTmroQ+rc8KZinnvfQR3ut5BTNHCZp
YHEg2VvBDEB2DVWb2tGqIvXQRom3aCh+zeCZk7h6McBW7FRjVNviNPGyiSBxT02ATLc0GiBVw9a3
nb/t25xx2PWAfvxkr2jnMv3b3t++axkp6D39yQO6Ut5BoH/xoQUfygii9vm9EUke7Y4X0etEsNrd
IjlSoQWZ2Fc0TnyDKAc7K8S2r9Op/B/1dd/m4Sbl441gWJFTV4RPpCXHI9rSg+YSo7R+rrSekuge
BuzsdskJ6HsP4ewLqoyw9SKn28dlGJVROqQrjk/50MzgWLUcEN2kCNtPvvYG8XcK3ueMTj8QF2qj
puF+RzWsUQ6ZoGGc/2FDTl10em7RGXjbf+veuvJgIvp1W3LwK9Ipt/8/0Py6Qz7MG7NE4YHWGg6S
ywU7uhwojjseo97/AJk4nHUU5VnFJhlzg67n44ctUOfajQUnwJFmCaeZ0Z9Eybc3c3+LTdungVjb
D4gvrPin2ejA3lQ+JiBSyQTG4a3ZS4EAsD8TPyZbeWQFxfAqYK8M5qYGkImxH7+EXrUzwj8PHvBw
HFe42V3XvfGoSo8sFeY6YOm5LYv4volXma7LGuWykatlvI8v7TJkKPG71xER9WjYjLVTW3aQnF+d
lhloBO7yAPDp9LzkdKhdddoqTp9LdrBp6N8ZnCPN4vKiTRuPioPsR18x9Xl31s4LJnr/kM+hxVej
o1yP30EK+XxfYXrCOOTnCgwAdCqkRfVcM3diujltoDaQK6N5Ld0FlW1Bab64yzklir9FzlJMDHtC
uaQiexJ+pMNUhv4OHZsXvxtw1w3xze314durJToDR5p+plSn6GkJskZKMAqz+fmllyCipjh+FKtK
JrK/Yy4fi51OyzU3mXg8X1uDNB8zJ8OUGSl4MjyC/rj1OLdb+NMVXWPeHbontV2Ayas0WmW/L77L
hB3LfCIdYJ/C/lgrAVCfs3gnE42z98E3SiI4LVleeYEWOW48zUD5MZnegyVjgb/vdY6scoec6NSJ
7cHv6hUX+B2s+TyeX0EnWcTfna9ctwgV1PpE5q13mNKIeyPuPgLK3W6GkGOjkIbOYdOSxNd049YF
tbZJozoG9ZAn7/VMRyspmef8OoqyFjsuD6mWP816cxLl7fNI0UCk/F2wYkIcYkj7dr1fnd3RtDlP
EQWz4Og+nRjd3p9QQAUQkk3gMIwVoVax+4w3PP4K2kLtA8BZu6mEdlW55ak4/R/nLeJhH03z6zsU
wn05L7w25TYj/iiB0qWnzrK6CbX4GV4VPqjsQ0NQ+gpN1an7EiNdRXUwzM8QFW8+ddyUFKsc2cSI
VaBh5RSZ1sDqzldg3stFaT1Nj+EkFL1BUxGb01dXXrhInZkDdLWkixGq+Fj832QbiuLc+IeavtTz
Ijt0udei2AJzHbvcTJYkN+XrV5pBmqKMI53qWircpea85Pp4gN0AuYIb1DQ9w3yKCLNuKPAV1oIP
cDyAwb/78UcIbZMYi22usp3ngexEH9K4DbpmZHdlCp7uEw++MqeGQQOl08KraRGITSD+9+zjdKcY
loIz1qzKIjGTrozmBGC2Dh6uD6QAeoTDOyNEw211hIDpgf9oUt+BQYky1mwRgkInJlqZwD2WwV7q
dpffMnYpybmnjQWCv7S1DbH5N+mocawYwETxXhNFQtSk3GwiHDA1YsQvZpzH1BkBbEQuR41mH5ty
ZVtgUVDyl27ZHC15g28Mxwqp7eNh8uybAY9wwA+gFtMPuoABSr1NKYi3c+0Cs+fH5jKJgfBpaKlG
X85K5Gmw1FTv23cOdcUj3yK4NhNZqxVo7tpAXG+fQ5d0mZM4N/NaRvIkHY2v0D6JhEZ/fooJguFK
wycv2w43pNv3QgvgWpCMK5Pr5XLQVv7MxvVq6O9AXd0qx4qm8cTXyswKrDP7jiS+Rg1WFiY74r7i
q8Y5ekWQSWdtqxDwXTO290eD3rSR/G0yT9uMOZdo2bYmOy6qLHIrjI67U8PTBPeQE/z7OZwi+pcf
kGJmdXzwe4096tOHojIVuhJAw+kf7Ek9G2JBsWdGnMz8ob/6D9Wn2eVzO63zDa+gwXnN5jXi3kRR
DtYbftg15ExnY7JRzEk/R/QlFfLGSo2CtLcbu6i6fW6iSsBH+f0eDDpVqNMwO3k/qsKV77pIub0G
SecJLtxLrL4HtowfUmj7IMJAGX9bB8jj23xO/JEhZoiQTYbgJEWwDvDJ7GQo3Jb957yxKZQYD2yK
lRRyOcsUB/BmiZODE4vmnjHoqCJCjj6htwKRliV1Kvz/bGGdG+72PjU9/r/udCwP3NTr2t5SSD6K
zPRlpCqpNVrTBC5Ete7Hp4NGFPT8RoJMomPsYn3Mbcn8g0XfvNv+HATITBPQ4JD1TxsaThXhsfAE
kyi/aG9NWxah6gnKMBo6rysTzPQ4C5k4TwkxOg+9UShKFeoJcIAkMS7CmyGyXYfgUW388UZKoFoW
rAilEYxkTG2+/NfHAMrBr8jBTfu1Nfb2S1M8qrsW8hLtejsdGeXlO0FduCbZqil5IQd/BK83ey7/
GRB94ENkko1hw8oQcqBUgKuvZ9pwR8vh0JNzO0NE2EFtmtMJaEKZRf+GQaPGXzCZyYRMAvWRBymv
bRGyO/1gJWHLEm+gO1H7wLj/fXUj02oX6vkNArbZY1393ammZjrWqQLF8wDt+u7CyTuyuJr9/rvn
WlHSIqZB3hyiFQds43dMj7RAFMZ+AZjhDu8K6o6dpQCPDxKqKJGPE8p31vSnMuI7AA7fXb9whDI3
UA/ZkCDZLES9g3V3gYi60BHvv0TpEgu62Rgu6XjGD2E3VEaWWnvIN/gW0UK03lldNJmQG7hqvpQ2
/8VHbTYAVp4zIuBrXXZ/YgrF1BnWp8/ZEnmxVCk1HEodU17gbB6hasufWprauqUWyfKI8ZaZl0wj
bTsFEpskBpoBp3eApae+JoXuN0L+tQkUCYQktpRhV+cyCbyAu+cy8Dmig8XQ5RqGnvKtR1RJ497i
pLuOQoacZRgR8GV8LDe7ZZyoxvU+ub2OAfByyq+UMh3XUEE+uL6O0pSyoMmozxmMY8pMsCY3rUAj
HvONfZltISuPV8ncqudonF28HoF2i3rE1cHYWjNthZcf59+4f5i0dffyIS/7BSQxLF7Ji0a9Ril6
KCnWepWcP137/JToI3mGiq3OhbrxYZg6fzJjQMFYPIDZ1ylI/NacYftr8qAw5fMkrhceYHn9OA4e
MhP2LPy6w0BWXBklRGXE0Fv01/+5GCrWsvzjr0VJIdpXMdfPW4lbp23/noRpybQMHyFW91FH5vgd
6421ZPEFQgoesjTylw+t/tpk/A+RipCYcaSyzY7TkDZrTeSZuPeAJFgqMcRAKGIWlabZiq9DQZQB
vKfID3zVg1RB/4c06xHlGzeeEBus5VnPPNEvVd8rYwtA7OBm128jLYSS7ngH4WcJnU9kTBPck9oT
2hP+AhATkfMD3hoL7uP2rU+A0skGEnPMTr6944kT5G2sw4U59f3IFY6vgkPjpcefKgSmmAktYxI5
QIhbJF8wiEWZ6AYiIRcQGFy7rr0Wm8uC0plUtYkUs5XBEvMh6CcRwm0ke5vVtzNNtq7KclIWe/he
00ynJSAewWCawvS7QGvQnp3IWBdyb6lxGfzIolK3wXTrobD3EoiDapRlrXDdNT7n+Kgo+oSBo0i+
txCMT5DJEAkmEuBzf0LJUP/81PfKt45bgqJRLTKCKL2mS+2VYt8uuceHAhWLXEuvzX2BK2DzXJxD
rUfcKlKLJh90zjIcU+AmBs/lUe3JS0mfgYT6JgoKZP2dzq1SPZpWJJOHn9tKYay872aYssrhcRDj
jYFTBmotHwMqvPWHRh4AR3GIJW5PCy6Q5nVxf3ViRiSPSfRl8SQ+ibm6rSQpAg93ZF+S3QYH2x+/
qaEm/in0UBIFagtXdquMkuo/TmWX+EXXsEzyOXFa/CiBtJcqzupAix4xv6Bg4zvkDoPTdQKIFeR9
jLTs/ZGPSwT7cHNU2coU2WIsOTc4TP0QOZfIx32VEu6jY+guZUXJLyBRsOxb7cHQvqvyUhpy5xDx
qBnTOt3vkNdxFfzl4oqH15e3svLI2E5TTBpFbN/+ZJN2fKE0MqLIdxJirTVJcVBa/sN4di5F0xXu
pwqAwssA3bHQiQ5ZcsXeViwTNuGe6qCL5QCzOBZ8YCWz2zY0/Oz6u7wtFqChL8A+Lm5ZXhz0N8cX
9i2IcsRSJtU/2oYx+85IaEJFK2Hm+S54RPlNG7YYXuH+uHFkvT7EFkDgPwL6m/7wtiataFk4XY9b
ndjF6UxT7PgieXMWfFeJj34TFD9UkZyyFqVrSgkhHufxnjlZ2vSi81Begyo8NifR++aK9OLcV89g
ASj4kxxrk+ayFzpWpvVTCZF0y84YhPZiFLyT3HD9kLGtWmGy+9e2T4fUloH+x2tCHlXC2Gh7UuI+
RJFD8Ty9rfbP6+oVnafstcQJegvLWMQzUtLydPOzTW1u7ikxUAncAXsvTv72NS45c7pU241H1GrL
uLjJDSygvEvhcHbnZABDv9w7RzUJklE+wRDwbZCUO/lcyBCC4U4P5+ttA9Copum+FqZ8h0aSzluH
vcBbzdkd0vyWkKQKPGtZ9ptAPBPz9GbpPivfKQum75HKFB4MFr/Y6QNx40CQl2CzvHop1pESJiu2
cBmXVABepS1YdJi+AUNB39nJ1lz2rY+leUtoOXNN4UzA6ZiKcnAZKYslCe3M7zVNg8Uk0yoPjJBd
EVRFmyuldai71RPiVu1hUYCaWsLpMiEcqUGX0MHpwbC5JgiKb6n9Ju/dNzqFbqryPHK09D/66Hfa
pH2aVVopB0EpMbgGhi26u/OGaEven23Ni8txhlnR8eYKH/UAzMjRejwMhgwTKr1632bEmPAIeTc3
fIHX0PIV+Q+FHMb6leXQdwWux2xxnseieey7E1tnf4p0QmCQDjcdLTVBcaPxwsBpyANdrKSVIn3j
53XRd0z1DjX3Herk4jo5G/EAq2pfik+UwdnRzUPsPPW9rmCHCZtwAh4GLuYOygDI7WvADHg2Piw+
pAosfpiIpswY6y/dHNI1Hh7OHanG0KrAcfw7SjghjVxuooPOc6dPwX6h7M4N30WcoFC75SdDkQcg
WZvuoXbF7C2emM2kXtaJqLkemVo5uX+pSI/KqAV0YBx+PE7yfwqo5s5904gmy8dWH3PKvi4Ms8vC
08kXdmJOxluZEuL3nJY9coSth7WxW8+rJWH8P46HZr+Or1XVL55qVrotyu+trpMEiMZHeFA0dy6b
a7gg5vVfe6ZsnoAbjQwbD+UbLhBWmICsJe+ZTIeK0hhvkcoLbzxkKBl17R8cOJCR7+pblVL+Gvrd
5IIKGl1DR83aA/7mDk2c6/Kb9DouwRPHt0al21DOXqyNGAyUoTVTXPspRaE7ahxmS2VkZO+QlBAr
co5BYqMurgR/0x/iu8MON5lhxgcS5TwxIpTzK7uczKcpxA8De72ndmHhk0UMjZlZJtsIi2JY81tE
6iy1YYF8oINoig4DC35lN4Ma9bY1WS28PxUIY4ZJUiu4f3ipNp9lY3Wknx8iabAj8dBveD/meOP2
xJi0nNNF5CUbe6nJkySXvfijyFBKvYWz/O2Jfz2E89My8dFTF8LFTpVHqDEhsoVrDEUMAStTuJWb
VoweYevGX6UIPXLGkPcr9VwRsowkA5AIZErIZIUmK9AuJbceFnpYDtGu9sp8pnE2Fr7hdIYbh/Yv
euC2hR7wovHjSiY/FNLuwbFWPG/P0nmkkDPPu9gf3uRzbo62s4cnEFZUjgd2k96fD0Q/0HptgrLX
zE9pU9Ntl+/nxFE3sJ1cSBsQTTOJqCGc3JltQYiZwDb7O8TDoyCf9tNGwP8MCW39/L9csVOoVbR6
AxpdkX9TTMGTQ7vUFB1bwnBmrPVgb24qY2aGKG05XTs2U8VIa0scPI9l6voDqtQuCI1BEZnARZdk
nWUbY4uY564FH2vDzeFj1J3V1wP9BNxCVPfD3SM2aRbKXLeD7cH6nwQBP/VzyCYbO35/lvXIr8Yg
pfv2GBUvAVKsjNp4UZLFBRELhx5yAE/yfnBYbRl+L6/R4y7TDag6YUat6+bq40fqLNqIE5QR2C4G
TNF9/5SFVCpaJ1tPeH3PlAAGLZsUJMYiZwStsinIfkDwTNvgcwv2xXBq2h+GBjF7kgbN6pAn8hT8
8N7CD7wdxC/1PzySouRfPvkuHIofAnETU6z4gK8RTez1EnGzXm5hL3WC47ydv6cjVZPAEinPUtm0
B9WCm/T+RP4oYzotMfUeKe5223rIiL4T72RR1bjpAvutOPzdFdlfPFGCyvBLXcYmE6Ye6+VQ65Um
snhFarJ9eQPlN4u3zFvgHhxA547UU9t7Wccm0oHoqYC3d/0ndXTOzgvdupYC7Abq+HXf64GnwGTI
KThIvpZsvJE0isKkYuM0MzA/X64uovv04kAVwmyj/uzpBTMx07VPlma/8nYnFGy2NkrAxAQ+rUPu
zhDLvQscFe7RB3raQFmJ2dTPjEdEn23iLbiDrkbOES8pTmDmhYXKX5QXNF5iqhQ4iTrp/nHyhEf6
dgUOp+gqDjxo4LafRjdBtxPZohqZauvGorCa4ugJxJUD2GZKRySUp+ucW2zftTg/SaTFJbcVqmHW
DhqQ8WggVBWpUHE5tEHX4n2Fcd5cUUOLKkVI2Ak39II8QqzYtZFTI1+0y6TqdSGKTZVngnyR/L0u
v0OgYPViNDBLC0/tPk8bWbz/+FoojSgRlNIawUnW6hCALPPP2/FIpccN0X58OaVKn4SZv9ixShAE
US8pfCEhYf1rHYvZWOjX9wgVYpMqPGVCnqP+0kdIJhBphRvtcaunmpfGM9RchR7Mys4ez70AvHaZ
ipFRReCrBK3AQ3kC47y8An8ByrG7UqKp3HxyoH3pk51TU+/AOpcuk9kUUfK8+zGb7Uk/ZXtpbQ24
58suX/8BtGW8fLQ1miN/9q47MKOeH02SYtAtFoK1Yw7a8vbG6Ik0kFgdimAHQGbG/pn+rqbyQb+C
hHcBICbzM6zx6IoIZLfe00/9FmSMLJeez6e7hvlx0SBExdA3KIFy0uVkWstdJqC18hM46FXMlWV/
UJUzka+r8o/nq23wKg+4pto52Q4RkxB5v24e2tsvZgbZLF0C6bbyJFTSDt0lfWw0cEplYifEiYpw
w26a94jV+dgKP5yJ3IU8A0edweydZDA0YPsblB8hO9nfW8xl3ZIbzVk/mq61vYspBrUY+jvqWzSZ
Uwhgouojy1oX60GOMMsTVvIca2+Of6U7PxlyWbhx9rlU6XCnzShzNExyVEkOSob+0ZhVXIAYg2pU
Y+DFqWQ5hvrtPLpP9NvSqhlKXi9cM/IZKJ4WU9hPfNC3s9e1DENfLUvI8M51vNO7anJg0TiFnez4
A3dV1DWzaOrT2p+SQAk5y8j9hDW9LSjfqrX2H913b9NBgsb32mvDYfS/MIn6DQ6odmtTrQFJbgzV
BTH/ncErFz4peQ5vOA/RzhRd+GtuHoYkOjvIh1CngE4MPMM2fpJ8LuHUsWkBX391LuJrTxY24Wu5
q/n7qaoT1Ys+/H5+VfrTXeG4V+3c9q6yXtWEok4q7dXvkoVDfulzmJkNPlozOni4Pnfqgn/5Ey1J
hpcB2G0WxbhJNQeH+Ns/zolxIK2A9f+w6MCz7FrSXdmkVJSSbXokLioIEws992NVF1WzDTKfEZLG
4xBpIlpVwm2r6IKuQBvzute5Zs20tXOC5qwkvDPC6ZfdW4U+qvQt8sURA52XUrnsyGL79lDWskcq
K0jIs8JEaxfauy59FzHYm1sZeeBvNcoiRTs4duFNN5NqdmujEfR0xet2TcKb7zGrE6U0cGZZEvXh
tWFtSjkFNouKw3NMneVM9oBEe1WEaoNZ1G0a3w6HJNdzQypafJlURxXwS1OXkK1vN7QINnFCWQUT
F/PRBTR0JJzgd1vDydupBEc/1lhnvDRizOARbwkjD0tsAoGXLbi0PLXVNQ5mC06yKcHVtCQLdef0
oONpUygQlhD5cunfErs/ADmnBkASGRH21pLkw7L4YqlwQ8RpSMuXLxo2QrSw0Q/q8Z69PjTJnM+F
mPX0Zg9VJvDoZP0x+Ltmqt8t/uA3qfvWHNrd4FxVe29O53W+V0+jsGt1IggvHLyzuij/GtOxotRG
cjJVgcFwF6F6udLPGTWCrV/y4fLc3oxvf0vVVzAKx+HnNeslZLXFAB2tCuNxWglb49xym32+DLbZ
ylwbWG2hD1DZZhkxlPV+a82JoH/7lvFLZv1J7Qfr6YPZN1ec4p2Ei1LDrZGcEKJpefME4vduvYz6
aH0EJKYaRVgjlUy+4pddQ9HmYX5yd7demhnMFLjH+WSdPNZSi82wED+Nb1AScc4PE9X7zd76gj0e
V+EddWwGVsD96ZQJvdn+fr9sodC2exfQK9Wq2BwgztKWlQUrFSQ9n1FIES/5hGL9A1LgC5asTDUu
LoJpMyP8EFQcl1QeG0lmZ0Orr16e0GIU7tQKDLrEiXYEwHqu+YBqS9hedgaOaZlKfXf4Znnl4nc2
m5ckn3ee7NXyTrEn4uMdqBswSWeDsemE1/CdO7b2p+G3ihGBkfIh8Hsbv0l95jKCbAzeW3KoBTL5
DZVZBMRI8tWNevn5CvqPIT38pIiUxt+i7NXP8GkiXKs31etphcAZo7JWVUAXsZDeTRE2MQb2Alp8
4hPr6AHz0Gac75g4dzA/Bs9wGZavFGYWm/ZT0MWFAPa4SWtBFkTWo52WS6dmN6nD20DyVTdauUNR
6oenX8DhzE5EVpbSgJGH0zYf1G05Okve+j86ox3oXFl9y5Y0mMYVrBDamUIovIL7TtTn9SgbLNij
ASn2A9IU76sjzi5DZlE9se3mAzkW1LOAeYYm+b4j9Ft4LzwvYAkSP3zx0qw6HRQbVyUtKV36lY9i
IJKyqN6mxe8VIliTD/CQIPSS9UijCcbT3kbawdhwth9LWYtWqGLkYBXmyAZqPERnGDAgKvnFLsUu
cvlLb0lUZYKpaLOwPDcj5TIyfUWQG3gapo+UZOpfPL5zfgqtrgLSPNVaqocx+24vi42TISmDJYV3
lb/JWsHpghz+IdhRqMVgCGqMl2iCWQsN17Xczslc8gZ8qV6zjGv+vu1meP9j8x82yzB+VB4hDmHE
5SOOQDBnCwD3cJoa3ou4aVCjGiz8KnYFAS+tlkWXHaNGJzDJzHop15Ur2pmg0fOqwOIdFt2/2qmb
k0mmLEUPZQCUFmrATMiqXxlhjgiTdRflV7WIDjESTI+UoZjDuxgJBXgVhcFfOf7f7ThKy9iV+GWc
KJx08mQzF2tHALFpD1cmVHtN3g9VsJNw4AK/GETuyNkJl01X8wlLRg/yr7waAbeFYX2HgTV1FEtQ
Dnu5j33vX5kO09EAppgHJEUinIZx7NZu3+hvueb43J3VTKhVNawuWpaKNhKpjJgPP7BqxF6t9/7F
LP+feLRIYyUO20al6kIzSpxKQFxsgeWuLifn11/XowY6JFB57xGGl/IxpWOY1RgDE3u8mq1/UcdH
O2FwpZc6O6PTyR7Z4spXt6Ad+sOS4GejQiLf4bW3kjWLhuAG7NQXtdoB0ccR8ishtuKDwyr++QIR
3uiNp+C3y1SuV7S4PaJqQGa/blpf2Xosno5aGOY22kDEq9GvuL5FvCMkTz5S9dBdyOXVkSPGnXZC
IVKNDJ/VyRHe75STITr6Q2Ug7ZAKDlVMHesejYnKEei/Muzg+YiHbNXR0/ya//iHMAp7gPiB0zKI
5Eqw9mLiejiNR/PZByf/60Pj/7Lb2tIE/fPOehtfLGymdjxwJdsdNAdrTWwN/UgaOEtm/0juGETc
whZtDeY+yuKxQRN+jkPf3g+3PH/1QnF3mckS2mjxWW7gR5cSLXcQBNleiaaAfum1aVgQMIAnK1uy
8S5lkjwdJggPBjmdDNa/kQIAkklZk3VMzNLDrCIJWiNtcv7JGGL9rgviIgND8K/8SWxpBel6Z4kH
Pugc5l77CLChb5aP0lZzsLNZoLbGhPDfewcsIoUokAjTiW/PYdll+kicnB4teeBNB4/SFgH2utEy
n6foIoZle6cKVu5UvZxiVAFNbe5HyelS88E+e8SZyahyZgn2p/VXCKS4MNhKMaMiHjs9g0o7NMoW
EhEoFgX3Nh56DGFDuXkjG8lfJLCGvD7TjTFJSQPq8oPbcl8Ym/SuUKYEsKINOEpzXUZZ3j2cY62N
RNLn+U84A+f9eqtbT2ivRIpX2u7cFm1nNZ6YnkzQEdJG8ZKG50ejcTLYoEqK8RzXTKeV7Yaoi+GC
WhNtnJ5R8ywHbcvz+GyqnUgUH7AYwdlGUe+dC9SB1sC+tXkUV3C3Bmaw8ZBaIo0o0gCrl2ZlIsDy
hM69wpOCTUrk3jKlFqwwPbvgIhXEKw1KzEX8HZOul0srlcH1GMexpRdfwQketcunfd5vZg+ks7/6
Z6m6kBZoNSvwoY3snRViOTUDBTmMbVwuC/+2DHvHOG9xBcv4fcRKtW74rU7b2wJbZmxhW6VjL+pK
gkL3JDKGvYQOks1nvG/Y5hCTIJ0irWjCxbxhuNz+uTEghHTNIW2UsWbgJO+3j/YBG2HF3V7wOIlM
NWsaumltpXWNfbywWdnYeU/SazXmokc/+ypUpWO88YIKk8TdAS6ztDcN8IueUJ79kzNBf/ojNBrR
rxckjwgd6V5lxvZVzNxmrvfv760/nqSbuKqPXbSttPqHHV/0NVvcMF2w18TLEBWSUGa3JZ/y/vp3
kqOr7t6PY2zfY7YUhAThBTeb2jyR+lezItWf8L6YRosfpnkZDW5NPrO7v/mmkOH3UuioruImxLpx
dHGLmVQ4418jpO2Smqft+9NSBqEw0oueiIVbyL3verPSOQ5o/4eAP75BUPmf7loZbu22JBF3XSRh
vqibpWxfQZwG66eSa6Yif/3NxKlE7qvPhaFRLpAqOzpPtgHfXkmBxVhoQl5fBJL4HPpuc7diklZJ
oybxQoV/nbeW8dZ3CkRpAqc5JF2aWkitDUpZrx3nZCYifAtN2apTfdUSsHgVEuLEFgv9r3C7Gq7K
FrWzHfytghe/exMHwf8U4Emsll6YiXPbhLTxyYgzt0U9PVnUtRJvM72/VICfkx2853JalbDi6lWQ
bqMstNH0eTsVy1+0HJG/Itmb9FfNs+49xNy2QIy/K42RIykyjfKrQ01BZ2sGbuLmUj5WLfM58gks
In7y2qlxXa5ss9qt25RwYWxtP6iGOeUahOGtEwy8RoNfbKhuhOTXUBkb6DeCWuYBwMxu1ZlIp8a6
WACQZQvHbOUk0772AiDl+N893/cTbCbRqHYkKryFGSGQZIDEWzMWQY8O6czqdJQreROUQfH8oyoP
aiW9ogTfqTsL4U5dDb1bbiTx1BoN72Yp72yPb5/57lNYEt79wAgDH+7/eL0Ual04K2jminwRSnnf
go+aUvxty6bQ3BCLVYqoUI0JJNT+gNGHbc7ppjre0fJOnlmYUC97fpYltw4VXibLDmmshh1u5ITE
GBqxA1Wj4jQi+t+G0QfIIl6GOM7vTg8w7XvpqDC9D2lCZ3riN5AuDkrIz+tcvvk596PMCdxJLNsA
cjKcuf03ov0Pvdn1I6CQ9+FzVZb9axJCduwwI1kg6ewieZToUBilD0FtNSrGrCh8DtT55uJMCcS1
pz3G1VZ7iQxyRiPBGqFPpYu3DxEOGWGqBWyMG9WlXD2dihKQXCsGX0E48Gcj44xTB1JXZDbs+i+k
+hk0O4qpG21Cw/YhVX1CeTv6vfCY4o9YLL7Mp/CNVjaS/0qZxUwslGqoTILZ3RgGLRBrvQurlG11
k3k9aad/fK4AuU8AigFvCzFJ8vkMVa2NYE8IZx66+TULKAoPBg7wRp/EIJGdjuQMyppI1ys43CYy
FHffaKI8YvKqqpgIONE/hV2z4YUH7b/PdNKy3gCqOhjeEhg0puQs5x4rIE4P9r2swEtoVi0RPI9M
uoB9K+MFpdcGVdVZrE15D/zN6t206cePQ6pgvmCmOeYN8u51zC7jh0lEwz5tC9XyByN8ICEyXT06
Aq2EadlV033hGgU2rSe2HYWgMEYmS/V9q473FP3NOfc0mka2drNJiNpzV18MltWlpcwXS0MaBRsd
hA9AFx+HYANI963RD8KP/FuIgnQe1ZWOgG9E+TIF2rK1fH72j2N9zZdRaozW0/QgfONBtYyKd42Y
T+S0dCjd49vpjo4DoZnfzKoT97I+DJKttE/VPzScqZE2ReaJF/Vd5sBoQ4o6AIGm815rd2eVVngJ
1sXK1am53f7k8qyiD8hhoxo+prZRGncLDGUiaapQHCrOH1DICsHhZ53eOZoBzrDV93FYZ9nX8Qgi
nv4HpMIPRs5ppT8fBbixbBqqJo4bMCBQ58fSKSb8p3uv6zgO3BovpvMToO72YCDRStG6pQTxC4uD
TIPD28U7GeHBpfAs+pDN/yCSpFDfdRZZ7466/GciKeswTPe9llJoNa1g+/OZnZe9Fp4IjSowJu2g
HFIWGfgFId4MPIhY972gUjYpTo9vqqvgUodu9OxYkg5Ws0MEA0MCdb5gsl53c+tDn6G82hQTN6ht
S/QCm5RVnooRjvvaBxsTxtv+lxw2fDyt/Sxda/PTTdD7YMFs8P5tl8HZWTOEcc1FRloO1pt6b/E9
2r6wROtKL++kR0umcG2TchZYzuGPuA4hLuH+FswYnG/iKPL4OFkOuUVRlBUFLqpcjhwxcUTDU2yX
PGIEVh1QkUuxI4IahDk5gPXBwhQwbqFjI+XDY2jxu7rihLuj7H8Js37wVA7J8Uw4SwtRsvgT3yjr
L28gzT8xwwA5/I8e1dfRtnQPLjr5biB8248sGoNuAl86s/0HJXYkZlJDubiG9I7DG2XH4MoxiWNK
8PjwMSHchCi7QOp/1egw9X24n4v62ERWQ4KqXfYxhFtGjbzT8q7KYZSV5QFXBlO5+40FnJl1CIiH
MyanraKft827+9s/OQki0MJptvH+Hn1Q/rlkQ9C5zAlDlrclvQO/PSoQwMicJpTEMbbFkcaN213l
FBuzQoXJZd95yUBP2Uuhn/Nr0w4xkilbWu6ZpIw9uhB2AAGrQCXFI94L/DpXbPm8Y4oHJQTeb7ui
6RvFp5TWIf041CEf0RIkBQoW7yzoZhZ2/7C6X0HeN1aXg8ZsVaxA4EtQXHMPJ+vZyplRSV919t6Y
l5QEwyu2tgw4OEwmno6Kz3folq7Q0EnmuVRyfHM4SNvSNEDiKL0gOLLbJ49kNrxCq4AWPomXE0Q3
Weo46UMplqFpLcw/VCei1XE9bjOPkdEEFaD6HMgIrX8hYR+QtLk0SGFcLSrvrDlZogsf86CZiVsQ
kaRs2zDqVtUKrMVvtB6CqyEEl074PZHVmsaK6hOzDvsGz7LhIWNpW0YcTbjK2woeIyrzAAycrIy4
sSW0FCJWStpHpdMo8e9nyHo26+8yu9FYbw5U5dwmZiyqGQA1dxTpcd3wF1T3vPzVIlppQY19YLh7
ZWgHFbD/Mt2nUm2OwwNxO5TTR8YzvvJTkv3gX4dhkyXgNyL28MX70l1Pu1YpnfNc1xuVP+ha/yKD
AEACEBC+0IgZDulVh9nSNgHPmwrrqc3v2K8Gu0FzacKMT4mdomV+DL2KZCweKaeeX6llYJ8LTCG5
waXMCruKkTsu7pc1Nu48pJfdFyWp0SnqmnJp13wpAl79saLjrhRgH/qtaywXUMuHBHiPDMN/TJZN
gmcdqW0iZo3GYH4HLebZNcfObCwWnqYEYpgKsarl6Bd1GUQxVjMNKDJOFmupyVSw6vyXbj9yj4k8
CZpmRZG6n1MWWDVXvIUle9s/APXOOcWQAjDw0fN0gDaQcp1vanDMOIwFuhsnB5f1qlHsDft5DK2g
rJmRpiAyniCeS1bHDSf+JCyPiJrDs2bKb8Gjtv2pxseoGn29t23Gs8vJ5uhoV70dRkQKUDRzIZzT
oPNu2gU1S/nK7ZrsdwftzKxCtGTB3i7+a7wjv7/doYjwB754qLhofD1T2sVo7UDMkkhNq4DjIjmB
jPW3/IU2TnBwd+9sYu1XRbup9jkUaDo93b7EVLbQczVaQNYn4G4fEBHt557oqD3wGhg2gdywF+rG
omdk/6e9U5kEm4g8UCbsn/WynOO60x34xxSzQyMnU3uov3rHusLrrIyQWiWs2REg176bDWlTIWgP
ih61Q+QtxqO0GDvqxw/KVBJHDf2UhLHHU3u4pizVjN4dFl39zyFzs7lMjSNW9zit26mIUp9vqaVU
hc23WGwRkN+hv0baYUB/bnQdqurTfbz4N+KvsVEnTdfEedCcRVfv4PcUKE6SbSTeB+qfrczhI7V/
H7Id4p+FLyKabOSJkk0R/qPIx0e15DbQw3ECwIjfnHBKaxWyZIuHj6LQrbfSKTLZjgL3Xa1VzMde
LQSSeEExtpw3f9fR4z+jM8dk2K2WlSbSq3ECkdIQdWO8bGbeoXzHmwmqfcITxp770tBs0nvycWML
/5Z/+AsStRx6pxfPWIYFOGevan1sZPp+YFzShwzLmmAEt3tIGsCH+IV6explhQGN+cP+sG5UuimA
J8zSZaYUcmZFEK+LusB61BsPcjzCq+nzI5sVVtiFta/Ewn1R8iZGDYEeLs9FBfUyK4Wh41h8v5lR
8YI5QnM36wv7lUBJsz0rzqLXZ9LzA/tcQUXN9zKk8LnX0fqMkYVfcSoSY0auZsj6/4ZTBnppVXYo
Px/nQaJ+aEHvL/Dt5KDMs1ajGPNzqm444Uy524pgd0GMZxx2KpeKVnerDiQVCMFAA6Q/qL6QztW2
wOl4+RPwCSHxN4G7GYmPG9LFXzhw2WNaZfYLVH6TIcpL77l59iJ1LFSwUBF1YspyDDEw3WNMKOw7
HyDHjy/DGdtvs75oxQiYkBmjlc52ibj5O+VGqdtvv9J3CP2PxBzC88QAlCw+Ww5X6Oo1m8X8Yf7E
6d9Pn69sh1lTthNmiX6NRfqiXsqVeLpcCVb258HYj5qFmYIXPApCmrxZSVSk57Sq5H5L9IsbYzoU
FC8ppeUtGO/XltlOs4PS8x0pUSbF9zNdu7co4B5NpfJj3xEf+Q1Cvl08iSZ3463yTkbQc/BTzrc/
cZUceb182GXMFDukLrFoHJ3DJ2N2v5jkGjy6z1c8EEgYIPzZREI/1GlgoMLGIzJTxFyGAasqUlcx
L4RyfKDs/8+GJdZ6iiSeKArlo4hbm1fdQfbyNlbxG+O6QDWzJCCzdbT1wmt+IVB5z4F1nER+ql63
pOCHoSVc6oKdOQ9LczbSfpvhoiigTjdJpe79lBzLQcR5qoF9wCwpMN5EEo6Pc2fPcCY75EU98any
s315l7/IBwnxI5DWkYUAvS1p/Fu6WsiylENJ8S39lEfIHGcNpl+OXLAK27BOJCS+/6qKEovKFP4C
F0aJX4zrHXiKAHguUEiuBxW+hOlLGLDpM3dr80SByarbW4C1ABcjhS33+0Vrqm79zhm1WZpcRVCx
o5x8qCDzjC3Nh6R1blfKfqnf3l4KJH97zfVeo3xcyHE0VyDQUOhycbUeCbcSEDBAWKMEtUA35sV3
UVgNb/UavmfWnxbygSdryiKjBHlfqmm7fBeXfjajXNc9Y5q5YT2KPGIfjrmWM3+bvmAAgrkxkIcv
vEfd5+YI4HnHjrIEsZQwAZyauhQlcBqii2Z77Kc08YWdpcoDaHa4HyvHBzygTIj0viQEOALcyMwZ
JfmyZe3U3duQjt79bEC7NwjGhKA+cgvUrUJPErCnlFT31DGPxB2HM0uxgNz+lVn2SAUbEyal23MT
MoIt5Ww6U5ApZ8bX3iqkkG6j1UuItw/vpyB0EU7W/QjP9zIFR4PNvFs5hvDaP3McMEteVZTPgOnC
Khid5Rhq0Dav72r9DKSw7dfniMXH765X3GbShyBYjKuE7HCLXwbMx53fB5Vkl4AqXWd4t1M7A8yu
NWYJIfa8R6wlfPpKFPta/YOC3lJIuvGqarCvb5ufMwvAFEI3Mwuhqi5eng2N2DB+km347j3QshF9
kG6HOBm27SoKzqIl8aM0opuhRoI3+gzjnEAQwgbQl882BwtYpoljVo7lyuEZZXUgekX60FN9v3Vc
wTDZRifG8azc7tezDHu15gSpPQxCyNTUcVx16DKih/5FD6Osml9YbvGby8wQVu/81pcKFyWpu8Lr
3yCjzjRQSUCm8yTjq2jfKM3tcmfib1RKqP28lzTBOwdMrEN5m50reOpt/GhUYF1umdqH4CDQbTLq
Z5zfqMO9u1VisBDbMUaT8NCaF81x/5PbxbruJDuXOY+QgkFA/fPSTmbPDjOE4cb4UrJGYQY3XTru
FtmHIkDVyY6F6E7wkHkLgx5Aadfm2Nsg/ox6hYbhe4ze5inDkRaNL160/qz2mdVDxT9W0NluOiSN
IwA3uNpsFbZV6vxtUjNDpS0lrD7NaXhICzJOBs6lQfYckLGeB7fQHmIPgX+q6G7nbi5/ty/RNtjl
8ZeqPRoIGSmvj+rBLVT3+gBvBU3oKmG1C1Q+4qJSmu0D9Ul0PtDdkARUV826yqmEpV2OMFe2ubzk
+Io/Df48jzZh6eR8p0J++30a4sON8kaPffT6fyVX3sRxisHkC2P35r4S5v5lI3Tt+e82VC/MoYCh
9ImO30yfjSK9A3xMniKtAnuF2h/0ZCsHAkfccYOwV6K2tk82YzCXvxQHvqvxqr66Psu7IpA4u8BH
Sm6xeytu9pN73iRZF9V881E1VRvdBd8C6Cc/6fVrRg9Kho+OPdBNroRIv39yDCWjJEB3T2vggyrE
g7+wFAam7nZxvsAVffGho9zNlpsGrJn6xkh7VtI1I9FIo3KiOLVGzKL8zvcwDheXBjNHfCjmotzQ
0/gbisVc60bOShC2fdGqm5ZKjdxXoWHjDCaeeIY/EX5KGPqnRbTP10FWuBEcwUz3H7j+ft2NZigp
gfKh2b/fyz5+GCPQzJeXXARsZS6bSQzv6fqSSzUIqNmg/F+DY0UjFKJfyzA0BNWjQiYi/93jVnkK
r4cKC2ya4t+mNFpf67FCFSvNCDNPL9i4dySTOqlSApstr9if2ZlOWztHiMzjgBwFvGRJkCSSGlM2
Hh9VhxxLSzcOO6w/Jq9QT6aEHnLI8iyh15uYf53yeE8W7XizX339UiyDoz3POhZFD9/jqlr6CkPN
VgIFzTwfpY1bG8qMh2u4BM4CuqaaPnISZPZd0zj3iDTgMRJKlQ2Kkd2rOWW2Ewbb1tkAU4MD2aAy
fcP8Ae9tFD+z6D/hB1GJfVwEe/rngUSzYINISFk+46ngAOy9TvvP6mRAfm2To0GuNLMBnoIUueF+
wkQt/rmguz2gmZyO69+LbW0Mnngmm4ZqQVvbsZbplKMq09Ipee3Jz81CnqfSIK71ljwZULsWmenw
/zEySsMA6jc6zrSslzlpcd32boRBugbEf7/ib+yuDOPbWqWXX4HfdZW0adrI7mECoZuP4WFBEWyH
srUnmvNfwl4OY4crBJAb1DStkcBYSAn3LwPweJwsvsH+FrJ+Sr1SMBmfeLE5lH0zVtLppqqEqHNn
w/B+vzP2F+9RTu9F4cI3YKYuPSMIeI7MnBc3qzVP4i0JInSGjGaPZcA993wiEY1o1ZXzo6ydRxft
1tsGrBKDI7Fty/QhK34U8wAA713PEC8jLx5Tp77c3pi+SnytgPH4MU0x+PPPuk33TktfrVbQ4/LQ
I+S/zyle2WbNZuQvN6C3rSdMdd1Nzgky70zJgn3P60PlC8dUwWWqdMN/AybUF2Fc0NYfADrtv1yq
WvyZXhxofuaPRt5pJ+IZApId+GPYz5mvt75IYfKOBu43tAihkKiFnBsvNyatYkTo/Bqdzc93dZgQ
6gljBxZJcyPZljAqjNtUSNqr/1YrygzahldGd/z+mDgUQ64xSWiOfMVAvqg9VXP+Md8c4wCofQWR
0dDlG3GL4718eBMtiW05uhEQ0oyK4mW+XgicEGby+3vy95NKVqnm5PysFaleCyf3qXoozrW+pzKy
xeYzMDxCO8esHE+PXJPaoosrNJZPuHTNr9v+qeIaMJ/l0EAhtT42ydJCP1iAfYB01cY6DqudvlaS
UgMaoRQSSAPXKzO7c5D8zeqsqmnul+reePxjbBcs0EMsDCbuTHdAdbrTniz0PSiscnGLLzDlXau1
Nqx/FAn1OgTz4VuJgQZXef3QGo4v7vsgnCHEhTnAt16C4Sh9bxPOQjr9poSL32AgGKzBLmDQovPO
1Vk8j36pht9u9gYvzxnePXzhbqgCXz0md2KwOrNC0tjgGMONNx5ogeF424cz89LKBOyCxU1HbSaM
e1shr+Fw18i3/ibDdQKS/+x0IM9j/MF5wqjlrRObJXGyV/utBy1zTQBOW1BkPpzsv8UdPnZwJ02j
++Nc7yFbjEegwwo6Hrz9Bs8aAlwkCJRh1kgw1cJqxL8Egh/MVj6h+1rr7J3pjHqSDHsVCR9by4kG
TEwwH+zv4rsYKFZyDDB5E7XXkHSN7NONINMlJroGdG9A0TbRAgzQeO7kgnlO2odEIeHKXVQ3prZA
sn9Alkj/EC6dz5UCVlJAUDn0Ek9dtXDdBLG1Wt9SiISs/NxhRWxZoNE+vxvKDZiB/ab5PP28cQKm
Ws5dkExxt8hcUuylmteLgISjPhsopLe9U6UU3PNnnpxYnbJ3iDya3Lo6OhUjdTUh9qVFwXZW0C9a
D+uN8ADZSeJ11MHG8THPtjNLAnxDPM0HLo6AEC8Kh2JvjwvOWvWI8sFU7JfUJ1eLWb+WgnB4Ju3b
7jEuM/2oF01jXNVNBqXmvdFHbYxZA8juciBBVksrRCsnEu6XtGoIdDyN4T5dk9AWIkL5nFEF9hIE
kuBSVfBHjRqB8IANr4L+HutmtAgFMdWpqJi4RyWyXFezMB2vsvtMTdiKiT+L45PRgVp25EWc3283
xdSuVr/CsLKHt8DVHSPS/wudGf4fWw3Dnx8Ia9mQoYN88aEur+OOmo+Z4CJPqs8i4jZk32z532UI
JkFQ196L8Pcqw/oKTL70NTNzqUrO5qPGwwPPNBLwy8DPi8fGSpxyE/FU5wtqkXkrCeSinnEtFvNY
F9L85akqFoyJnOjPtRbLSaoANAOUAW5izOea8QNEgrHSoBt9ImP23b9rQ5J4/gy7+Run4WYeWROa
aeKYfDJiJca0eFwMJ5V1whhdaLnDxC3PytGlIIpZXKd7eDLpThyfB9sfhelZuDpFmt690eM0yNSt
jAtEqdV/snM7KZjoJmJQ9wsmEsKDaDCOaFydvxdV0EPoUIU3ApNS8c9QiAr0rmAkVFhDrFEnzqSG
DbS7BN/8OR1EFfjsQBDS9Mjot5DLBmSjr0BHidiOmO+e/E0dFIJZSBPEfufGZFhq/FuehQgICpHY
naCBKeCMQ3jk3GJr4dEyY1p0HLz9wHyfQQDw4FYZRM/Y7NXTBu25W4xMcQ+2mp+yLz34uZujvjEV
KEYyTXzCJ6Io6mbltbIdaC9lCU7DWfzWHtHLU/TBO/1nO2bgRAd2JthoKAWxMKBrhcSNAH0wegls
PT+QevVeBs2kEt6k0FVrRVb+v3fuURtI4nWF/FNG8T8mXvVx7E4ouGDYtfO3nlCQT6XjO765vTL4
d6cHL1BDMgt1phhsI6WQkTa/sb4ASn37ao3CKrW30XTz2WH4um1q2OMBOw78U2WFWBCRmDGQq7oM
23i2PI9vEd7rx188AxDUkZY0VHXrCNH2VFOIE9EG9wBqHQNRMeGqzU9knEowmjHr1rH4sOJvXX1D
48mAx0TBuzdNdF8K9Gi+4Vpn7VKtl0SQhO2CzT0U2C/ooFxqEqooTxfNke9ZxGDRrZltVuiBSJhW
+IpcSDOZpEhRngwRuiJZKwAXM2bIyW++CoMSGyODsw4j0QR7DIQ+rp3CvyWhmbgSzMX2Jpn8lgDA
UTYn0fA2/lKuPVV1nQyJi4AbHfILXHgRsfz5V8i18OrCTlvhImcElUpTMTLSPTe6uvUywrlsSFKE
7DDqvGafgztVgucdZc2bJpTPqn6OIerItEs4ZH9Ai2xLKm/tlc9DGWlEA9jxRag8DF18IS448Z2T
2YuBMuw8i+d4zem4o7ScrP05I7RMhKo/48mPE6sHJJQapEhWEyeHKgVesNSAHx3ZTqezjFvEtfIL
+5Ogsy59K/K0fL2ccKg7skOuA43+QC9OZoIrdeH5sUv8OZEmphp59MqAQONs3jATXnuS4ReFTJKP
NkTFcoukePLC9v0qcxGggKLasHAOCm1Kpvt8a/bsy6Zt2dW77Zsw69grSMg+BIPexBwsPDMBX13u
uq6kjcUI12olyhzn88hB5vVdhrx7Oc71zLGwKe4Ln1fFnkdlt/6lJsaa/RfDfshqN1P980xBVxB5
HynU+IZ6+nsu9ypK6uQz7928vFKnHNvI9+9r9SgeHchdcT3IGZTzvHyUipHjZ2IjOhizrG01yiuB
4FkgjnMcNNLHF5vg8WR849v6T/rUKNVzDaERUl+IyVVDGDbVGhtrjmrLbOC1eZfVvV/hR3dr1Tnz
BfTW1Hg886kiDidrt05x+bfAzCazC3JclYlaavtPByjbotggC1W8ynGC/AFxHG6BtMDpODYs9uJv
ai9W6QaJb7XV6BPPQSSmLYfPNIX2JOe9BY6F/JiropFnPaLA4Fq1O6Bc4fFemmCTCeTcYZR3ZyQI
xL0D402DXGMANdN2gUnPFCZ0KZSMTgIKqfkGOR2wS7F1GDDZVQQa61EYedPCcevLIGrZEQieTQs9
qQyDiFlMQ5qo4adG1cT7in/aybg9GuivGmNc4P4dITAgMPlC4Z46d2JKGAkZs0xevlt+PFevXFZ3
C7xJb1C+06tPbKoqVDc+u8ycF/N1GADJcINp7TSCL4p1r8IQzZ81d8WshuWSZo5SPvQTuZZWoUwR
PTKLqNPdKYySjnODd22s+8fXdQeLNUNzifkJhUhty197cUUkRvQ0nvOETQ+rcI9l3Rb8m3oUe4JG
rKGyoEJBLyh70mlAuIM1GyeZlwgmBj5WWoNANKTiHJmZtmOeK3WQaPNVf1F2T1355VAivUl0vIrz
ujj1nh563chEwMkANfs1UKPCw8nXGRhTPW2gAzFwt25+g8+FXDeNIS5izwrWiDVlLL7RwnWCzL22
jvPKUO6gQO2gz7wntFInDUk2IVm5sjf89UDBQ8rgU5uTqzewoL/sPqj8FfEQM9T8ZZF88MNNf2ik
i3PsspmgFrj5Ef7e7cEFo2qAvb0sD0WkHX8V4pYoVtRDuzh+e8TOgWsJoTuWb/LBrton0CDYM41N
wLwMksk3KOz0KJ5+l+cb/BPRiA18xDC0/CG6qgCP3X2O5oL8OhZxc4GDxrfoi3OFIQgrCBNQz1aP
Q5xrV8kB2UhP1yi+n2ODge6mfi/Y1yTt1VdWz/QKOpRE7Q6rJxrOz/H2MJJnZo865KnFCvBgpRrD
jdF1O/ZeoZhN37sQR9MsEcIwBtuh7yCP0mNXmX3O8v8lxz6WKwB7BiyH+b0l3W4m8uxXVnsgZOWA
ZwiUiVhjuSQ1lwYCfDZlt+C9WrM+Wy40CA588PUH/6w9mHUxukukL33dQwFrDn3OplwToVunZply
20zHFTTRSMns9KaNfz6rLaQamdE5XWY5T4u0mlWH+VSK+2WBrL3ivhvts/L3fIXGkh71cGcXua2K
v87fR0LAlQ+xBLkUsvGmEYCtFDKXWGStMUhnwOg9qNLP23dPrVl5kna297HTxRsxnEWC/R4Qmcln
TB09CNUFUxF8Xr49yDDCK+bjR7FGNq/A0aZh09rKHAnoTA0uSqOhMJbcC60D4x+AJyMFyCsRy0Qz
AbD2AiOVALConcTQRRtO+9h2yR95bzCYvP+FHCpJgIBVxa64yOAjNbz8+UPhQKtPMXJ1PhIb9QAX
7lp+hLr37txNNUxSp+Aw2ftdWtaHxnft2/rNCtYcDzFFlUkkZHTvqd6JfcwL/VkF4VXxFWlXuIhi
pAYM3h3CiLLL9puWZLiwjQQtuJzYqwQnhcdcy3HaJw1xfRlLI9iaB2LM3WPlDA6NeI6i+5lm08v+
LAs82jdj+qRkJDbwaODz3k5yec7nahsXiIiUFwChwKneK46YzRS4EK09r4j5iuLN+A7AtA8O4d7l
NQloFrUkZiV0n1r4kbDtsoYG1H+CBTmiuu9a1Punxp78lsq82xxm0BQf1ykcIczN2z6Yxoj5J2Lg
0V9xg9ujcbVN2XobM+9oKIWowAHRaiorrHOWMO8FQD5JYtfOQ2Jsx2FYuqbLQlpXC85xcBH32ni5
lPAtGvvBVd3iyTVLp88DyxIHg6LluK2J2Tw3yaEGZHQ/uxiNWJWtGK4eLji1DaDyBDJg+5uUPHhW
v/ZwHie9tntIgcobHvOuvWTxNh9hwp1pMnppJNhwWVbIOTOM+yL3Q4pm3+SIaW6jMKlOLbV+3ASu
12tH3ndkMVCEc8TNLRy3jWeHXG3qTpDTrH93zhM+jkR+XtnvggNYUJeevr/DD4wPqFx+niWdhd25
bpBC9yA1MjPU5wo6nB/pcDEw3c4iqwWtZEx8Ef3wt2l/ffpkRF2V7z+YhYgH0XhIF9/MICWi/vox
uzSRtjbXkfXEunS8hb6ZHVF434ePqgkz0VGkdu5sSymrdab+YZN1cgTFFmq3hkNtg6+KtiiszhsS
WFPx/iOC+du2fz1gr0VI9IY/IR2tk8svB3BBarERp6KPiZLcPFwtrdwzm9sTqme9jyAE2VPjmPw8
dRDEU5x8cv29wO8C8Ab1Q9NyfEVm//RO37erEXNHMRGfO+koCTFVzdpXkfdv+7CIclZXtDzZHWNO
uDtwFLT9UCxmxyglYnb74j0fdl0l7Iey8BegNgrMyJiS8EmGY35DuKxPbj3kNtO0iYWdQPgP/cO0
XQ647DdKWV8tP+YLU/0r7xXmj+G9ifsjlUJ6EnAsKesQeTf00o0nRlrTTfzReA5JYPUabhq21Vfz
103FZ0q0QnKN6fuxlq1J7IC96DLIj0/766BdN95LltTmMSxkEcFioP9scp3oQulyibw8Uer08ANL
CPSv41QgUkL3ju98T642QZx3GOp9S4d2nZvf23sakBvNQPpFELxDCaZVmlubgrOxL9nRVz4d9i+u
P5oUSlRMFvP+xfimlsJaDGwn7yE13KU5krHAdVknvvzre/OYUllT4z3lw/mF58fcr3359+9kn7o9
IgsVJ3Y8SluT5b5+KiYP8FwgZogCkYN2zJAeJNn098KtO5TRl28AS2WeSBO7OIZeFa176X5k2H//
TrKAvWfbDZOG2Y8cMjpIjUQ55T2T2zxw19XlyKkj0DTbdzLDqM7WzLg9MfgfUHZEomvOtckbq30m
TID7tYZf7AReDay7xiloIZWjwXk4nMMsu2Da3pepIU2+mqdvzSVZyFg4yuXdbBQoEkvVxWdMZaQs
FkwIUpzqewwRuuTY2TpwTEwGZVkZIdXJz1RSRWhAXsHXVh7H2St3OPm/YMgR70gz/PhHr0oxBecT
qKyHS3tY6AB3+ucpB60t6jL/Duo3+lHNBRNsVka6QeVRCxpmEE3b6Nibgh/spiNPuvF7ze84QJvT
+YKAJLvJBN9pPQGAo+PK8eDoSBypAOKEf0mI0RY0dQFluV9KbnJmLTUrnYrfi0bTfEvTkT/vA0f+
fR8ntXtD6ZiLpSAteIHowqX053p7O8fmlNH9EH5Gr4oFpHSxTHRVCVzV01DfmMcySdDgkyzW8GH3
L3lI351oe3p0XRCZeiC54voejW/CjIzTTwRL5z4BUmI1Qd7v5yBZvbrMT+d/+4QfldySpsQzBf4R
mPM0dwQk9AGMdFpo1ixY8ef/FtOsnIv8DNphoU6F0DVpOJ0dr/v20qBPOWnnGlU7L2g5LR4v/c/E
fBjel70VONPS3NlV2M+2l9vhBYOebx+Uq5LPA/9T/iKBgA8u0gW+xZtDkjDA33zqkR6oTDxWmMyk
UXxqHLW5Wc2sesYPifG/j/pwSAEqjqQfy8SPjM3tp5L1r+O0mii/fs248cfpf1PqF0tddN7tqbJM
nAFEbQjrgnNoVZDLgY8nqs2lctu49aK6YZGtqQI8nzG6D9qMtqb/J+kTVtdhDzVmfKYT4+Nnc+Yl
SJw1DGCciz1V1+m64tEkatNAwXRKXMH20fC7WrmN3FbRg+p+izKpe09xDptfadfC4XlH9L+79PK3
CKj0YuHb9/Z+8DUFjBlH6QpV5umgv7fr2G15GfXWis5AmakYG/ugCE3AcvBp5tMy9GHNe3jh43BB
lRt46ma8LgBaF+NgE17+VmIO7w7x7Z7wLTv8yhvYRqgueMzXJC4S5iBZ6/rB0Fg0KZw3BuEGOdSI
TOkUxRY8s8o8qHFvtMpl/48H1Wk8RSibwRSPDVk/iyVgp963i5zOj79G6CtSDxVnrXnkZKoKeqaI
dedu7iD7VM/nzSapwoUz0spc+nYbqBCp2DdoeUdc9CJ6xoyIjkW03FC6E5m93uyRGddX2VkR9m+p
k6QwVUp1zae4T4DVMHC8vw9EV4b8IZajmfTqkxhas7L5f8D2cCX6+m1nkBaHNoNpts8eN6sUlQMr
dCJknh3MMBY7kGzMyUM3sdJ9+gXt50D16uprfkXzVE3qUwDZU5wVeW7X+5099MCBJr397zC/I97Q
yyys4M7Eib2S+vh1VGlZCAuN+nvtDQhgH1gTwcfxunH2UMY7bNYFWnMVt8QnfWd92QmPwn7yGZ8H
PF2TV4WdovC+5S/9LefeI+brD8X+N6GU9JxuPU8Nu1WwKXY7SZvAeev1zVtPrvv04e6FFgv0FaNC
INn7J4E8gnMpcJipGepSY1O+KNgUnBdI0+xu2p7NztkpPvk+zVhnIBQ7eJWJtK/dFQpFtTW5kuMA
XBJ720oXon1OF7iH9H5pkzFaKjbSQscN4J4Z+iciVeWb5w90dlexx9HFGICNdKk9xXXRjX/QE/0R
9p1jxUHjp7xI8mYhlhG69EwjvgUe5ElG7DWu6y7mfBbReQWvUYfYRwZe9hpyYTUQhxjDuCwilgqW
ATHUrxQ4vmbEsXpbd+ucLQNAvXfV3WJMDnuMVE3Gm87mZ08vngCNEAonw5aB1BNf/FNRzc+WLq4j
1nApjYXWMi3itw42uJiFr9qAgRjaWBzdHv63Cf7DWsVgBTaJ21OFvYGmPnW6oZyKOe8YcqiIuJ6F
K9yHvX2SNP6N6aSbMBd+XN0ik30BepYkZDxUvitei8jSQIjLrEnU77A9t0CwWz8MRUqJUhYxOyV8
tmw2woDcX/jCUUsxqyrdzXU3c6RULFk94vsZGkMPtU05xK+ZkKTh9H6K/PZDr8N9vHu632mLid/u
JVvILnWKI83LcLzH3390SOLdKEyYP1X/vPXX3B93Pog5bOR6AVvtxIB94bwPGkG/6g46GF/BCvyt
pv3UNRwM6gR7CtqlSt+1V+Tk+87aBCaDx4eZwQCggBBIklYZthdofQIg1KCNeeOfR4mYEx5P4Xnc
CAW/QwI+xFiBGye2DoikZ1WAQkpfzmntVmXRhlTHAyOQq8P57mM16WlC63wGPyYuSDlyvkZhOoOV
SBSaeF9p2s8Vk7r02d8GXSZao69nNLDaou3AoP3IK/2gfP6FPuIJszAjiRsRVODBmwtczT0FeyBN
USAzojSKcwhwR0CG08z+U0lJjIzFpSW8VfjQCdh7s5ensDpUgIOncdDLumGm4eJ7kQ3KoDyQloTw
YX2cqwBU2eUZnPqOzlFrpt8xkgp1lq+Rr4EWCD7tmqSCPRIpEQAsH+22UPU+MYbY7pmfiJ95D2yR
KAER8+WpgxQ/pugrgl7hXNh6Q1Lsfxx8Xp1jOb8Uft0/wGTBSVttWtBYpTZ8TCoZ/MXSJQE1HPzl
+FJdxLLz2akKB3UZXO/jNrdKo82YZc+9QcXWr/i6Jzprom0r7x/p92eWLMZD/ILbNrGPf0WRgbzy
pEFnTg+sLVAdCiPvkEWF8q7bJrKOcfmOTN8Fq3aoAaPcyrjvC0v7OdPMqx9UOBzzRZiUVuqR8A1J
fBpOn6s8ngNw3bn9Zc+bHNndUtwJv1ptv5prroTKG8SoVyeYLGvPqlngyfeQ4jzOKl5lgEfxBx/Q
SS5AskdJs/mcfSSNVg0OOh8Pz5YUnlGmHA2zk6aGscyvzIo0Yt6YgG2nndTspWTcBB6RTJh7tsum
GvHl4iSxeDYkM38kwvE3kppuE24xHlvUe9fb/pnGN1W1GguIEpv8XtI6l22jxy3XYXw+AFifFgXu
FM8hQxLkLUoMzIUxDBsad+Kvb5C1VMyUYrk3vE0u4vVT6LcA2bxbnzg2HJhe6zfcKYn591ZwAbNt
n8s9dyLpSg7Dw2LYRg9vEMa7LGWFI7uldcd8LlDmSfh8acjlb2QWHyeyNFmOBzjO5kDrEVEtd1L+
uSH51s3BRuUPF06Le+tzhc+beRkVueSmwd0ATlpK7BqG0N9l45HGGU/BVkFsW48PYvPaF5p3PdSP
LFtFgff5Ca1i/mlakFRWuCuQTrNUZIln7G1Xr27B2TqpZjVwP4ptQKzR3GFEF84z77TZPcdaVlyD
UmReARZipDYGI2bFi9CcXuRqM3mHpS4HBDtjk5NngDnX6txxmNFekFF0oBPdCfeW4BiiS0V8naWm
IFlPlY/MQkDhv12T9yRfS5ACDkCIvPVNkJCsn1KnjDWNGTVDjAe47YWUjlQwVlS6Tyl4GdivxGE4
mkUcWNwdAUXi7kQm9SilkwEEngs2Zt7H4Epc1q1JRoqiUdf+vHQPqlJOxL4uiAGKxcKVEYzr8Tnf
bgudONNY1YtWUpyrD9SEH8xpIt2uwldwvSMWWBbYIs6F3xrg/db2I/gME0fR184NJY+Fl64Bv0XM
oz8l1Mh8q/ToDbrEyV4nv3s/Dj1XOp2Zk7+Lo3OL07cic6FcXi5hjYVTugBYVmW0cZNjyfGAlFH4
sOcbTbvpIgrqF4iZU1pmClRcOUF/S6fXF6zvT55RTMG8fTjenO93bCmroS05CTafr/3fjBnbkPdF
YUyXmPWp8VPvOW11GwvhI4yjR8AKB+C1bAW5SC8aTkUJ9wa6j5GCp+6qe1A7IlHDVpXd6xq4FC5h
LfCsE/tKFPwwbZcJtnEGSxROAganFV9OL3059jdkEHSj/h4LS6kelqzflgfbWuxPu2RDwoBwrmC8
5QF4PDCL0m6GUuDPeTfgil8D5naLi7eVm10ZHbvm6yArau8u2PsreE/6A14VRh7L9+t37vmQPfPE
g0w2/WcLNn7itGMOLPPDFDwrbta49ZQ54HoSvnTwbrfnU1EeDVrRjvpwU5Blu8gChshOHjlK3/VQ
brWhcIef/ml+BNyhjlbOG7gyRtN+woI4oYfb7DIV6SIAyyr5jT2ko8XBi5V9RusDBvAc+OtRxPh1
G7IkrKCvR1nc8ZwVe3P12FxAQyA1zUZhB+uDF5IP+w79pxeZUVP/eICJIFsdZFNDZgQTL/eP2m06
hKJJq97xP+5kCf3KKCsujmXqu3u+3fOA6NPCIF+qMme7BVA/lMg5hQNxhalknuzMJaDGPWhAXUSA
rvsLTap2KSDIw1m/3xFt9jpbHN7dbTYxMsJxnh1wCBsGn2Wq7abuSXFGETkwT6RZWIdCCpihYZHg
kmXTqvpvtiXBP/vDcK/lV+RPQwIonKQIPcvwG2/4vc0ty17IaqCTD46dELlVZX5Pxm4Te4cB4aZy
mNg1R13uiwilw4HiRCcQ1z4abUpFXWCCoxEznqscv9Ko4qYQCvfDwFnBHvMZvGQWWCDQPgVYT3xo
INemCIDikuyUdnBMBzpN4rUY3CGhagZ4+7xOdhpTshBoGS0PF3qkbB4IdndkRMpa/+lHSV3qWrKC
KDM522GodL2d3bfzW1a/DDgURjVUhHs+ZtuXnEaRGFVoypzjpqRK2PH75s2U3uRi2W93ubD42S0t
KKBXYUX8Z2osqQMaHc1BCVMrv6EZ3XOxdP+DWMSZ4T9RCM7YR3WFVGXXKdw6mb69vIvsZVt58nAH
Z9ZYivep3iTjxklD5bwVDLktkLN/9+4m7Z6LEbvoB1G5cmDwIIvsUrS2FBs9L7V4NwzUkOR4//Of
KD1tAQ191rFSTHmwi4RYPWA9f2E0F5ECeFXGWrvBpb5zliwBQ2O3bSTmY64f0aPgr0aj1aMavojS
1B72venLBuSuY0R9kxLvae+zsgp0gJ8iOAB0yMubUvRzphA6L2xok5cZg8Vr+cTYQsKzbrUY3AA9
Bggalqxgh4D2YU9CitRm6Xk2qugqATphJKMYR1/aklvqLRSdzrMFevH5qnAi6hJJOJHT7fs9pI9/
S9f8lhmEyPaBFf4VdZvSogqVlGIrM1dWIFAzjUmm3XhVdG2fWtPS2FEayEssxOGELR2kP93Lw23L
L4W/YEC/ukSBN+D62kpvcaXX6zaq1zRY3Ttngn53lEq4VvLi9zTfcqY7yiRktjz3CtaDdBYNL1xU
9KUhOjQj0kS50Sx2cHEyfEPtFWglxEBvtE+hP+avmwGREN84q5tIaCRgA8jETUBlk0V25ft97jzQ
v5XCFw6GY8naZ3dYnUgC/aXZPpcpi11tE9lkW7ysLOoPrVRfNlCk9M1AbmQ6cff5rCG78Te0YR4J
/1rdAVIErk3Y9hoyvcLh3R+r+rpW5WBC5mpgX3bGessiZlsNyO/Yc4D62AGmT6qPjaq30LoSXalD
iIU6SMGZY2CjfJNBCMTLO3+fGgwf06f9O0ifvbOG8chmOXps/eHrudGAyhmo65rexaim+2VLLEHG
/Uveo6hSE5n/WQxubM/z0C4nEi5EYPQImQJccNXdHqGa59Wk77/a5vt7qi03RQNecmnLCsF6HM7A
HSsSl+McrdPPH3B9r4yW/MSkesqsG7Pv06RwrB4QNiHacJuT4Qk1TEpian8wxytl4TdfDRxESNGs
RDzZSiTOibSYCcOxqFinxwVt9yFbDW7MIfdd6/YHjL13zVqtlvVlb+/UO7Vu53vZy/yLrJKMYj8c
6/4w2jMfutRlnmaV07wE1JMC81IyL4InkG4BZOKTF+L2+Xz/ucaw0Upl+AHDLOlAMRWN9vAHQc2E
W8cOPJT2iJyYQF7t2jHrTo/B/zGhGZTL0PhYyaoqUJuRjOSxC9tjYc9Wbs8wUT7V0n83jkCNNAju
/Tw3OBserO0b8MS0Ab5lTBSAxXkYirZ9hex/ewmViyYEH5/ow5S+FZqXd/t4FG4TWbZn5zCMNp3E
QQZQI1dWT/ljRy9ofKALyT3+m6bljhAs7LbsC5L8t1x397fwu16FFzLPZt0xfox/9jMUE10Z389l
chen8kbjWhMhAvYPfm2bAqKCQu6xdVgiMjqO4MYCBaNDTp8vWHUGNGdKhP1RPkQMji0WLvLVbja6
RP4A4RLc39WHtWxTYPbHgNvpQruakbb+2CZFLJ69f9jQ0WmiB6wx+ooGXErBkNbNCPt5+7FRs4Er
Q474TAAVey9z6/jn7/ivMvydM2xvqH5KsCIqRYLr7jk36+pu8BrBcK/s2JvMZX2dcqveaPfWQuN+
Q5fnoL9WUGrokXvdv/TNuSMk/tKFpy3HzceRyPzwdN/IsFVWBtOM+NdLJTAyWfBdlKAzDS/ktgqG
VkqCSxjQL/5EX/acwgpoSptbOsN0s6mPkGXgc/hfIa/GGFFrZKygAJ3R04h+/UC8hCz5YhMkZC3g
b2/360AfZANPUc+MfcQGj7j552cMx1rVKR/iy7piBSf/i0jbHQ+a/TzwUFOwHLfnEr5WF+lI9CDS
/aqkAEeOijWLZM57B5Z0QXcGZoYRkQF0KeJ2/DSxz72fh2KAaZ7DCGB5PEHWL1HlxDwRrG5ZSi+o
hcasDca9W2b22kB+cCY1b9yEv25/5WwDENleQiojaPXi41woiJ+fMcrrOpeKHl4Q0sSCTRsjPYrP
APvOdqj0WU4/CI/kuTI/VnXKokjpHaOYlymnEcPsc7IYdWhiIiSZoWnbIJlRKPLZjO5m8+6ZTwLd
PP8g4ejJvebAF9O/CwoeKvv2/LlFYxxulpOo76m0O90yz0vFl8CVp87XFJ9gT+YqWIxqqc/Ik8Md
zbwwPY6yRk/uFmw7t5oV6E+LRxaHWPliapQPwIAJ5sV0zuM1QoV1stXZYRsycPBRq9jS0oxuCEq8
S3CU7lLkn0KH/RKu6MWS+lWGCsO24Q2iNXZEc0iScpD40Gc6ty+HPFUxwfW9vvwvmbRG5kyqQlce
f/WPn7pXR/He9B/L7vVusM48v8ucnE9m7sOC1Nm1cW6cPfBx1dvsgmH80CWRwqblXeWarbalYM/f
o7/HDQQUZDh0e7iBRAMFWk1F1zKYzVh47ZStyOsBuoNRbTY9XJ39SC1FVkSIBMAc7oegqE6nhyR/
76yLLeVFy8xKSkyD09ISL6wU12xwoZfeRVULG4hvD/yHVEPRYJ/4uhUh82bYTV8xzFUyOvpuTVAk
Jqo4HZV9r0iA61K22mKEBhTZSSVGeS+NqnSR9zKI7riWeDSRKvqxdJxqbxA8+oIxth2oM7vpiowA
88usrtMf9Eeg2LVZiLZOFm3/JZL+hYvba3Mz7R2SpxehxDewfcuOQm3dfal2k0lFA7YsU3bBC71B
sIwoS9qXs78OlS+14ULmojI2QoMrx9nTBC7SwN7eQmunO0AjcHLOo2CbxX5LD+GXfBOrXRGhggG5
/MnjOTk7gl7uYnTeQUjovJiM0vWjje54YFCiu9wd5yaAYJPK84mxpWshjXliSLeZwAz5/T0U2j8a
4S8eDso0+zQxk1F4n69vR7TeudrQx9D5XRmOhTVI0WNyMNSSkgISM8p9Yzu47foU+I3onutmb4b5
lUXpc7MYjhtEyHUKXZNTQW1qhcwkBGgJvnx3tGgoDK5UWap4E7oq242c1B7c8f8bCP3W83yrPPKL
4fuGHR3RVDNL7Y1WJgbBveoK9P0ueD1e6/XhppZfBiKTKpJ7bm+mp5AjsgfGzpYdKqLOvtmavL9u
0oB8zqsFA6XLNITE4rYowuZ+ZmBmphTtmJ5fBxs+15dnPR9mAgHeYvYy93kOFuvHO/P5qM5pvvay
HTnxtoDoHCJxbpjrlqUbEhmCiw8iJpMJ6Z3mOuaXzrxgkM/Mfq0msfw5mUW2gN89Bly4lHeotTs1
ZSZcGF5Eh++o3PBOr3W46e7x4knHAOtFJDuiy5zbB3Tf7PXauoV83a9//zSv+cyysqpXZl+0SVkF
JJKaKJ0oWpx3CIZ/Fz3Aag/C9ShFCYzBWDpKGBVdbg8MXA8ikTnC+HqXhklQoricoSEXmN3lEwjf
r/E6cwEZp7QJREiJP+nY/6JGX2OT4XWLqx8PXGdkknEbQkjzHzyYteSce4/dIRZ5eDQvw/UH0YIC
BlhGWzM/6TnLVzT1Cxu7+0gmKM2jvjRJSXIGPd+6CvckmqC8lDxCKwFWo48YZ8HrYcmmRNnwogBB
B+K/skAvgREJLX275L19HQSYVGwr3LnJoEvw1eo50jjS6NPbXUTlE2QFBKUWjP4pro4ffKkyOYle
OkJcC+VKFaBxqSTurC+WhqvssDqQacQPIVWsAPofv2qzAF4f14c5oB1DdB83FyA5hsXzLao1KOfg
2wtzdBJS30Lzt4jkjRBgLJCWHSh+8862cnTTrxxAJbvKN/34+cvgWigR3Lq2PEoH+sMct+44uVKb
Gd9moay+PDWoFL+R+QBKyXfO57Du+1y7GyZX1vz7txAddAE1ibZlUAQ5ffD07RzaWhcfhHwXeHec
lZxBV21wRrbeHteb18zysoHp/WRNr3WSkBdOg7FjJhMe5Mk4VltMC/frGOUJECDsK4d77bB4Yd+0
bLYfx4HyiiyX0LsKgmaLKZYwZxED5vMSow/egNM7QMfsfwjGrjmdc8vNjZ1BjCNPcSvxK+TghyUx
4aCIRJ6dQdj0qLgCw7x7G+nvtt8Ckpj9axuEACGpPg8N7rwiweJvOxjq2ealUiP3gBRLMyqKc93k
44FU0hwx0WNHc7JxeqWQUunsqKvRY4U1fPtsw6tAa7uneuqTHa5wVsTw3rCzOdbAxwHGMuaNKw7x
3wDobC1HxAXycD5aTEZxHfMowTp404G2FLJdzadJQUVBPCUHktd3hIfEZkG4fpOzZw0UHZQCj9rS
5JuUsD9wt9lzA9A3oFFbHYXSmFkTHzo99CPoXoS0wnjYitHtXpiedzSEytvkNw+DZuARZ922J2jK
tKLPqUqRloe19u5z8qOYbpSsnWVQIP60RTXL6cmPFCLFu7/3npy+Kw4pqO6P/q11m4emUMHZ2vuT
fl5iAD0dmiiel61Ko3tKExMmOJUCiGiPR4U/TMV+Kt4Tj3scVAP/jFxojjVFTCTw91Kmz5fGw2HI
cUQodrieuPTUwezm2RF9HW5TsqlL6DiABVloCYGoOuAs7UaOhj2tFWXYV4FWN5Z6v6rXbKsaXojV
N0hAkdPFfYXYh0o0nnnPZi6zZcHwmpGTfYyaCL3LnGT1l/qswiHXGy4MGiBLPcmakf4dTb/4O9cQ
iEnNGNikQqduF+K0b1KWhBWiE2Oaxkx2XIH/oYhnvbJ7W6ZdCnjZuVXBJMUYmq+aeBnma4H8pZe9
rwAr+gMKs+yV8xRUz/+1fNSymPD4Qs7pDgFW3Q1YW8p4PRKp+Uv0X/gbRd7VnQRdWbe0rHr3RFMl
wMQj4JkSrVyZ1mwJIbao15FDkzKOQs9XcZOxtupjLBAqEZtOxDyCeItyfVMkfuoDXLfsjsHqiePH
XyakoXGAy+UqCWkc2hEK81SbuXxrTOmjv7dAfVPAsRCLyO8mRfqbd/2UjR3+G1KRQZwF8kTy989v
BlGHKxtbA+u67mHAs1aKmIKh25sCoy+6OF/gZXZzqqJ8wAC3ydxQ6lWKKOoMeQ3f7Q4X0srRp+t6
qKgeiWU1WRzGEV1IogWhlaLmrPqrYH+m1MNVVuUx6K6up+2u9APTyuLW53Xcdht0KMlYpBd+cKTs
AnIzCFwALdXB0cGeurIxzyckTDM1uuzYQdZicIXdqgLLlAUhwYFYIczaT1A6AWTpV/45yWjbwQYp
Y+uKHYv9iI+ECv9orjf1y3D/0cFXHQDbc46C/cfoWfHhcjjedwuYsBsKbGv4BXYiJD8JX0SJPcWN
XtlMKJzbKyxwJhS7jy/LYTRINjqYrItE7qn7hTv7LyDP65tsdQuOkEF85Lp+VRbBf69Z4P0mgZi/
cd7gbSkcIPuocyAVs9kcFM8gWvgtSGhLatjZEm4UmwgT5DARTqcM2EiGCEV/1I+InBYF2HtrjDSt
YIfRtWm338awbifSrd921pykYtZidzNUSXyw4aYdTXCFn1gh5FJoo6oN1LFHBf0u78oIZ7yntFU7
Cprg9b1C/cwUblBACyMrEl5Df7SzgDWFQzV9zSz4vkD1hNLlL79DFSPjqsRJDDN1LR/BGYfLRD5q
pSDBAlHy7OP55i0br39YkZubmwiSGfs0l9tQJoXu8FjFsutbdtUiYR9bJFIY4gvNoRWPNo09pJ9J
3KKgxRiUPCiERg+d68Yc/UTGqiUxrYbdSE4E6W2gcgrDYpAG+6anU9SmuXTvpFHnAdWxiNFK1+ad
2cEcqkMg40eIS+QxQ7Y6/XeKvlHQBaZQBmEH6wIh+3ibwlyJM2WKygXy1zIgMQG3Q2DhAwJM5N2D
cub6sIY9s9okPu2IIpEOVWWPnm7FH8M6HA/OwbhVOvO7iXyq760Nzt2YhLaHBLIPeohJWD5vWfeU
IvuALCngeVAIM0/G8sH3E3JYpS25okfThX7QDi8KoBqB4snT0leuWb+vfjrKMRQfiwU3uhHqEZys
YrSmn6hYtNQIA+bEzKNWp6L6tkBzogRDCP5Q57TjCTLt7ivwz3D2mx25aS/IIbUhU5d/lFnUDr0P
ZJ3jW29bfzswTWL/zO7oEDQ73lULLY4zP8WfbsR9bCb82+/lFry+uXblyeL082sgdWAJTwQoS0gA
Y0t/E7xfarzxZBVYhd+1PGcC+R0wdcdr9uCAFk/6UeQs8eTfRYOiwQfwFJi8hmAvU4HU6S/79rc3
zSCskKEvN4dbJbEaOQcSbkChZOPJO4qXaekRsvuDbJGzxwBdtjJMKXwKekPUNoI8Lwn9b0/rFdUG
d5tIIN+oAUYx6+aLk0ShHwQLetbJBWK7utVv991mzlDpgs832o1oQHtPbdXg+jzV+oj/JHcU2W5x
yvaC8upPU8q8CI9QDZaK/5yeQLYXlzNxTfoPznrpWyq4IGPjggwm9BSMjUEhKB7SunOxBzR8nl0n
WFtyqOdn1+TOxltGauAuBC0YeU+Uhnh7w0kp+XbxgSywGeNH1pqspoXtmb3VQzND40ygMdwEpnjN
oox982Yw992RqtAYpsKksCS2XPMVxKk/BiCBg3c7nX+mU3w7gfitrhRvx8/r5PBkUgLeCCdd1QzJ
brJ5FSUcAgh57X25zwKlMwphiCldN+5UaU5OjWCW/2Xx6vjJOSv0tCTkWTGzN77b/FIh4O+zp38S
7uAdCqo5BmSPpWTdk3vaWYBScKn4kJym2149IPNyIQxQtU4zaVEFNt0YFAonwIw/soo7lHYG6izC
+neghj7++SplCVzOqhcwJvXnBQ4hlpH7lMQMNdL80Ayj0Lc9Wsm+6GWixTnwD2D2rMrY4I77LYHw
IOe7XcYjNqCoNLq/hzyp/ojybAHiWMzbpJyP4/bEaVMBbgYrsBaMv3qWSn1X/3gUsYiZlNPNCQh2
VkzGtmMEeExxChz/jiondlSkP6/VlWwOcs2vuZzf6weiP6hTKReP07PlOQPbbgR6qZPKN/EvzB1P
vd+psocVlQHnwkv2z7IZ6gmrd9fMlXBk9+/ze2jDjgkPC3WjVkCQ3Yz3pZHXp1NoRlZi0FBWLHaN
RK8OzEXPTLe4UeXNB+0nEBv7x5YgG3TB4bvbDluapmcSWTvQl1IJsImjUul0D87wsH7cPaI1aMTO
xaLHp2noMBLo+huN595T6vIxRbtawLiYxspDZSgCM+wSEtOWuG5vdr0DpYI8AQ7BFLkB5nl3qE4A
2ZJkIO+RjC8IH8vNX7vGIbVxKwtXFguXIgUgXZJR5xPar5+a/2xfmBOyBXdnBLA6JvxkleQwjlVK
IYmwYrZGXuQCrBpf5e2eZQDW0Fnmegek3WzPDfffLDOWQ7u8X5x6amndszUNGic4/pCxvCpiVm8e
TUzkt2EYabQ4qWbQ8BNE4FfiPGBGvWpfbzlsY5NZ9X9X8tgcRA96ngEbbjNBeWtBaeslUmYKKU62
oHBeiykQXaM7PRinHXoKgzOjVqLNafSPenYJEiNPrWnrfSymC4GDymnHzcw7tt6L4gv4OanYnKuM
4Y8TJFNhFOlBS1DnZMs12G1NvXn+JUyMsIOGpPBgTzsW0ai3/+9jpd/ssZv6AQUzBG24qEAZJWLA
zY2H78caBSo9+MtKkXkaS/8WKt6UOte9r91bMhcY8ULZIA4OO49F04vgwOv6/kRckBMruoHaKRFa
tLeS5tA3VvKijfY2Z2H5oN59NJPsR+YOBJLXjT7KZdemS32QBKDYPQAGewTMnDzOXbFe5MxtYfgp
L5LttxqA007HK+W+TQKobC1juAeQY8SJ1837vfJ70eqWHtiguTEmSStRjUZrOVr9yI4LIC557QoI
I+O8ilFTugpPRTeor82IbMVFrLVE7bPktQMUERsZu1EhSXM5Pi3B5Tl3mW0uRpGRFpvHZCweDjVo
2lDYbcfiJSIrZBS0HDtsvQWDN1hLKw5SZYvNbHM3dtHLqR03eBnkWfrEXMzi0sjOhRjcSRJUc0dn
2BqGdOBXQK8aU2Qr0YdwV6kfzlNiIu/PtCyF3s03J2wxefGBK/D2QBeUMH4Dr5WdothGWWrZPncp
Cfek/9WrLUMKXUm45I5q+IKJTyauNkrfoLdBaHVEOOLNDSP/C6Evss7aDr+Gep+MW70CBqflBBZp
kvwkGNV+ktaA0mu/68ovGEcPf2jYoyAk+GMfu8KBS/tl4oIblksDI4z8YBEXM6U96xwUMd92gumw
veQEYH8rAJkj+L1GzLHbMuSlJ1ccMJl6kCYJi3j+az4eS/QyVLAcbK1RIjENXUV1OlbGW42o1H0W
JHuOV59e5FpCZm3c66kB1TYx6fPAg0BCdPltoKfjFlVPr4LMSW9ln9u5Q8dG1EX1XguGn4TH0KLb
Rqtd+xrllYgIsf1NcVUA+9Pmzaj3SLGI4pJoASrdzv3kV+RIp4EnLX+2K0ETDcKPXJUWycdNC2SF
Iz3dq29d6O1LWjfvniK9QoqoPlNQSBePJCJuIpyKaiILy+ag8L/wx89ITUx6lgG6aputGUDXRi1o
06D+RiE3tjNgnISkjj3A95gU8G+E2EkT8qhdLwEsdHcLyHBo2Hjh2VkfKHqaL6v29u1A0BsAj+N7
D4tzUq0ERhheZ0GSIxCNcCfxjsKZNMlQrejUXscTatcH1DjuLGkxKfeR1eawr+hoNMwfTYcruJE5
kKSqEYwy1qWw3BdhXnEYvw9Sy9IHdCG7GQBvkAtuU3Q+0XHlpo9flECZdD6/kddadlgXi39dUEiZ
b6nV9Q4QexA14hfc/CY/wTRdufRH0ejsmaFcB6adoNpt0+ypuhTdeOGnaruD+sZp9TWxbmh0MhtB
h9ZEGpnTyySJTuGWbt8f6Vzl3e5xleKnJ+Mw3Nqrp6tgfzpuTV1Up2M+JR9rnkHwUbXp/Hzo2OEU
BqyjqHo5r45hdp4fkv+vvhyHcpeXrMe5pIbyho6XxNbqR7IL/Vy+3jwjYphUmKtTInyrENanjJyQ
bmfercInqRI0g3OYOrfLkmB1CE0sMIagwMZceAzrIeFkHb1888sqa7cjn/pmb923ZUedgfDCcJJs
3E87rzNKuQsn5aFOP4/sw0Cq0FobSWke22mPPL9NLAhIsOBjLMeqpZ0WOm8HZSzlLGdzt8oQrpsa
zQiE15RMm6VbkQzQxr10q9nczesi88UiyJQY14yDI6BerK/iHFCTSa/Q1feXXmosdgBw+wmWGb9x
pVfimioyQ4fcErEIG7FF1khizdLLDcBUjpUTsK/tBh2XbnOJCPtmLNZXV6lWIcIaFpes8YUEgvv9
M42sosGms3+6z96xqbUgwsRqkOTvC2hcIhKa8GKs8287aURL35Xry+Ha7WAkRcRNOVYU7xjqdH95
WxYD3BXE94cuu4LUAkjOlYmHW6PsZHBCPfC0kEPEDeg5uw2/ElSiPPBxAyEubWtL4g/6famyyJ9G
hvFA+WL3dVGmkvWBI3pys8QUul8RhzFMfi2QF5tAj2CmmAUFi6Vp6KdxnLti48AeCh0YPPrQjKoD
bgrBgoN9Dxi280ev+3gGN3GDbH2wIenjHEH2QSqaTOJimZF1dIY+OTliOAYeJrqDIPUnOndck17h
20QxhgRZlptVhJQFwy0XqIQIunJTYv4DoAOlpOQiProlBVqxgecKyfv3AN4Ru0/6jyBq1rmP93Uz
sHLrUFo83Z3n0wx3Gt5CTepQc+4KMwfPx5ZTbDChNiB/SYEuouutiWeqHuYYbAD+r0AeUvg2VtW/
nA4OGqP0T9KlN/w/RAHSWbKUV7d4vVlmTucAZUGMsZd3Ga4me3Zdmn9I+wUpcvKbyaZQD9P6NAKg
0yZ2G/qIVdCOLpnnwKCNGfZV/85UIGZhrwVuZYYDhtIyt0MpLw2o2KfqnjOwyIFjNc3j5qAi1KwN
JAULd2RjGmbDbe1a9mXFUBUnZYqYdapKMqb9ytGG8fOuVRcWtIHRQ5zycNgpCTi2etkp1w8x6eOV
dFW0cW3pgZnviEoTSVObvy5sysJ3ufo1n353yeci6PkZ6ruZcIjfeJYhuf6zWa436CCeqE31Lf+G
Snpl4fMyf4pNYLQDlfE6bt1GbMiCUcgDII1Nr+LWNZLZ7ZtxCqwv57P+yR+HgsTscpCnQ95CCsJt
QqeXBb2VcAU5+3u2mA+EJaXmXw0NbsDpjbFvLBao1l3Ksf+0gj8MGrCEKFaYHU0GkZZzphRwIUZl
4dAmttPxymIhZtDDBDUnAMcezA+Qeot4CHFacbEB0dmKIxZBaCT2J13oMhoZ0/B0+knqCMlrMuHH
IRKakdTenjxt2YUOzaMAMm8D1d/8joxjmWaX1Uf5PhZ+psQ+6JaNtfrguhWyxB/g3jgiKiw36vWZ
qNZMfNtVj5qCCV9G/3wx5QcCjTRaVsOv8thalddK/MwaQdylcGerXKgYycEqT5RmcBifVO8S1gCI
jiu6e7QOFrHvVjugsElFYYxn35zbBSyEoiUiYWGrdO2bpJfPe57tLphIGH/4ap5DzTJmhaiB6HOj
kLzmPeCd/324pqDwBd3ujTorMZHaN2dRE7NA8xGPDsr9cbO3MfkK2tbQpwSg28OXV/LDZI3lVlRE
rdba2QTp0qV1cHPUCIhCWyQW6zYgXaf0KnmMCiZ3Kjle8ltqNc1oteVBq3boPhy+OzB690NpbyBx
49pvGLhQ2Q79xQPMKnZ8IdOsEk6XD/3hNTB+PykZstTiO72/99UTY2sQjsrQ7m1eky1BJPoFMzSg
4DPINl53FbFUCHEvXf/6sQdIB5AnzJMKUjJINs5gU5Q9e810zZZY/K1A+XDmt2OTKWpXlXOzhX7z
fV9pK0Acl1WUE2+HUt76HAHf1MFI6WF+BeAUQ6qITtf3glyFWIsaJozBfVnlCAkU8VisauyCK6bv
XAVOFtc2hZoC8AxbRzJPGf9VVLN3bbYNAasEUGeX/ErBMtNGHohQCuCYgJqBH/geb7I4iVpgItRJ
dvq1JhA2m9X+AMXUuA8AfOVc92tWZipn8/RKdUS8xUE/ev8q9ADsc+JJSSksCqwUg7qlHZX2AVP5
1o2UHyKcGfXBGlaDq4nuVw9q0Z6vaSlTqRLiRjlT1T/18nd4ay8pxlGjvIvBsYpg4q2U5aQg87VH
/0H3FOP6j2JleqH5hvrQZmK38Vv8G0A9GBX/nDCAE2ZLuR4ut1KaJayp03+PdX9ctDXZRZ7kQCiO
7gJirduU5h3NJvtzxdsAaIxHCTbPAagKtgBHLkFLdWpJYINyYK4Q+mUWRC9YYOGppUfNpmuqEbyH
8LoC+oqbNos68yq+hWhRd7MWJI2zjYvoDkjOpE8kIeMlpWxUq8o7xCH3L1HFByAXy8xCean7MDDn
UhuQrL0nxvweG5ZHY448hX7pctWtPB57wVTTjakhsTmlckUaqPATCz3ibv8m5lzGWiwCu+bqnaXM
s3Lv1Yewiffof/Nams2zSlBeaFJDjra29l3fMa1sPLZ2cCdzqf4meRZgu/ffVhJfTrvtdTxbEMJ+
gJtHxw2ngMSNzb2cbbyCLNVn9qssQbelhdDylbh0YxmkKGgLNRGVLOfpPfJq3snrsbhES6D/eKzR
XzW36IQz8j+wfP27v+854WcbQlX9OeBH+K7LurOJEcYIXFRCBIJU2XZsFZrbe2Gg0xdDUH91gjYW
h9i4Ki52Q/2taLpViOVcXGPwKRc8EurneymWkrN321NlmOshlsJhUwCaYL+mDyZIZQxqhKZXmht9
PUs/GTOlk2j7zu1HSnJoXEouraZK/sixWFBZcNCkvC2SWPgDyfEdT+zhcclenxHiwVjPSPuqxR1e
McC1ihjTjkvTkfrjcDqlkg4iXUT3XhYm88xoa6TpzjmEtNQXTaGgpWxJeJXCxdfMsEsAMqS/BQiQ
AXVxTwo4MtY/sqm6SFIgBFMw/2nlLhS+OihHyqMrJKZxYJD3Q6pPxGI3jiwMeAAr6eXBQd8Q8c0r
n6ASelGy2R7/mSfgw906IbPQ4vGFWhBryCCHHQJ4BrEzNbtZ40NMwyKi3C3Psev7NhCV8eddKHif
BXJKKAsC8cI5LYOsx1bEhD+Z2alEELsVsAxrKAE/rz+GaTOdbeAVA6v62i5FskRU3P5dQmY9mjFZ
TJkFa7+2tqHwH5/kqKdS42WI3qe2gzmkOEcO61RGlRQe8/SAz5vGo4EI6b6bL0JsIQQstECeBrds
gmvy80cBbeunZQHdoPDMf9ZR8SUvqJeebfednoATEcNUAiELunBTzPyFF0C/15pIIXmi4qXUbyiW
ikx+InOdruhRNNUde3fZ8kHBKUkPwTKYp8aMZ3AoGVr5eCJUH2igTRyjTxtY4/C/APDcoZySOVpx
5FPffgr3ixa0vRqCoaYlBm8x1aQG964vKptvmC4231Yj/9NESI1zsCkewgky82VnM9r4xiuhSlRF
IOiki1R5kXPW0w5+u038u/BFvq561/WGOPGVn0IBfPAV0tdDd5nvYz/FrOhs3Z/uVLdrST5/MG07
qcky3xuaNNEdCzyz+3kZhcnryV6kV7TimEjMBUFqDzB8u8QA1+XBgd22n/xBbkqJ9hJLvNJTgDms
i036Nyb9tWDpSae76vrCPam4rSkdn4YZTBZ8Yd+0Q2i2bvtVSin5gB1YHaRZkBhGAS6OmhRvMlZz
y3FxWyYP1ybZ0Q0VT/d7Ju2Ayu7YbuT5h0aIvU9N9KSF4KCBfUf/c917L0To+ryM+0hrp22412dL
9siZfBir3fSi0jnSU1VlWBFJ6YceJ50b6x5YEBfBGl+yp/tCQMeK1YCALu8UiHbsopcVrmRzW/gu
HNe9gGV2bN1gxCjA2d4wEGeVn1uWRaTTNUrrxwneg91AwIie0n4OjZqwkxpbu6OFhmpZdFbTa+a6
ib/u+f8HIWOqVPeKYUsiQtW81Lr6qaKtkOzZ6dLgK573nHJoMAdf7OmL8zI0tz8mMrqZMzVKC/u9
ThAoA8/69ukxDdBiMrOI80b7NXILKP7grI5/33zybK1beAlgpKOiVopS63O/OTZMGUpcmLzHavrO
hFeACC21EE63aKWjIgCxQPBYFz5aJ5wvmq7YTeqoTsF3YYkx3mC50K3PBGo4t7OdKbdR30YqTCm5
YltWIgSmdOM+sKpCXQ2/CwAiHCcyHmpms7nYm0oFWIg32T7rzq7w2SNvOa53Ty9ti19Gy//kuz70
3wI4HJwIN2+oPzni4u7hdTxKLxooYCBwQvyqFMijK2dmkFlLQAAR7AX0PyOnBFxFN09heZpQuH7Y
VSm1VfdtPGf+yWe4guE3NVcUKaNFgnMmtLxH+R6Rk3AFdJQ7c10czNLvFUHa3rvS2NlKyi4JwiN2
3bHmr8JVDiIxAM6GF5aukgtIVEw4y7oQxZqn6EcC2mE8hgqPsH2zmX8vrRAJV5fL8YRBJGvRMcip
5DL8khW5yoSF181917bFysc/3Zx63+ptGzDZIp65nGYrbJFkgnQiCCNF3QqA+Vi9OGVSx98G+NQw
qM1H9LCxpOIZduIPebJPrtHEEJUzNgrWW1ZH9/Kx0Q/dKaVlqvYINAkkpDY+vU9reKEErZX554Kg
m6dgIHowIVZiBTg/LZNeU2b/IJ5lInP3AETpxCK/i9V48WjvJ32cQ/9q/yoefIGW6p9tuD98rTCq
lxZoIHHefPrZCeK11PsIQsuM7TQdIbNFnWY0b/881j4ed3qbXLiCjVfg1y/rg1aF5HhSTjE0qK3W
bef8g4V35HtrpyvWyY6zhBkHk8tLUEgDoDZAX1+825E+Bi4oP9X4EX+4z8pdsuXRJup+3F5g81/c
4rI1Jr60+jiJR98J8HCQW8LNpgMRK14N0lHa7/j6VOUtAvgBwnniXklPtDIy4aTiKfB2MNTd6wxJ
A1P1LeG4/SZydGDZTDWbQx8bQUmMQApe2WNcNnU0Sg/N2ZQ5ShtCPgzzGH82Ev06lPxGP/rpm/8u
RdMnLahhs2GBAEqCmN9efIwz724C8feo6M+dHVR70sksDMocM7WqbEiiKIIcO4JZ4jXtCAqnlGFF
oRhJ6rI1Ue4w3VDdZ+dx5DmlhAdlhAt8kGsxz4FOBW8RM4Hre4Gz1MviAlZFFvBQxJNtbslJjUbm
O2Tv4kAy3itVIE1/415aGjTI1aaX9nZBDgOcG9ZTBHZyE6Iyoj41TM7qKaWlgZFRDOBr8tuJl1e0
zTcRqmx0Mu1QruvfGRDiHd0CISuVfYWvDcgm4wVjkIMoWWNu3FNzZd37nYeuvD8xXKw+CbsxHMdF
jLiHoXJ6SCQHW/vwPVjxl4dTOqP5IgbeQTR7Y7x6HldZgPmTl82bOcE8VL0aht+CNm9aZait3bnu
3r54AfbsMHjymUhnGRufViI0WRzE3bk5rtBUrltKPjMvQxT8csjUnk4d0EMLvTlzfka49ax6ha8t
iLg2dYJ/88w+qJIUww5/kgNTRUQrtApKq5FH7QbB/0OTniV8Bg1C/YjKV3DZumqUTC/O+hZQoltn
DdwZy5RxuCjMu6d3WcvxeWDGmN/Iz7fXqXglhJZRwTwdINzNvute3h+4vaF+fp6ju1zli4xN+tWa
DcAxn579IAIUvEf5SlsNEP4LfQXzdoUnUycm2Ne257oLi5+CWOb3Zmc9ODrfXfSpRVgUUs3yjiHk
dPSyDn54JYqUy6WLEcAtXPRC+XeS+fICu4ugP5evvWb0tB0/Gv0cU6d+k5yHfV8B5PpKg5n/L0zw
MUp4lY6mIFucqgX5kcAJt87TAwwLcPpojBO5tRCqzHJTnsfgHAl9RtV1F167UJUjaQXqTf5eDmOv
k28NLz5Mp0Xmgo9LpKM1L8Uj2gztcODWB8WX3+xFj93LfwI0owKwKH5U0ykIflVKBEiSnv52RnC4
yiMVYcN2gnZL/T05V1eYhI8cj/WUjdvWuRxZo0RIXd1D5MddPjDEo66nIUwmEBbsRRsmvnF2SUKR
EtBK+wMzh9Jdexye3j6SkXb9KQdUJG9y6Mo61vS7vh5f60OivKPigwyXrmXFjEDzQjOitRPWQREZ
jkXA3QA8gHFZhecdT2O9ccMVnmnQzJrufDKJ9KJf0K0ZZFnSg736BnNToZRMjYGE6X8ee/VFQYr/
ydrEgAVxNkHPXT+GA3M4Cr4QLGa6zTEL4AHh54YVh7lNKSm6bXJCcjfpHJbqdusQHg4GpAtR5pZ1
Em0afFrtjhrs8U1x+QwFSlR0LXR/MyARQpeuG2Amfo3o2jOAdThRGP9b0SHftJn2Th56c3+9mzRc
2aDL4Pr2KDZM0G3I+yrF4dPyC+TVDIvgNGiiHSJ+AIJKruu7T29bhhI4OP9aek5h21GfAouAUewv
Y3zZ8HJ5wgp73Pl/cv0ckKcLN3h8yGmAiw87qHQOix4uaXdlE03430eOiqRXjIKI6O5ivTCGTH0h
7+R2rPdbiFvTnKm6Q5seRy0xPG4qyRCf6dzo9mQ5S+a7t92otupPwGEVNjlosJmq1k2xHCwdmkzf
OmLfYecbcTWP+E1GRTnVxzOT1uO3xUIeyXThfxAXega+/D3jZtx8fTv0eI8z3BbTobaS6bZpOI2U
Z0HECpNkHUpAQ/YBbnSUjcsCBr4HHfM8bb8oAJE0AG/qvCR7wX/Nr9IdDZHeK6AULZzxPHWDfNTk
qftsM+PnyxLNC5oOxt+snAtu6FNT6m44OLTQwKOqL7KYzekRVDGCuQ3iAlFnU2m9br2N2n3rFwdX
s8MCReD+68BnVmcUJevQtOn4ZEYsJuKfybyUsvDKTbD3QsOPchdxDp31KAHvHiIWeM2UTeuT5y17
FZhWfuq5dUqz05ullPbj/+bR6MUZIMYISk40+5NA5lSaOnSsjs2uMH/ozmirjATiezymsX69aQy0
Nw6y3fZnXWK5F12QOUVT6Fcgx4Y1OYJ/bmGe6mooBma6uVMEO5VPev+W81b7yClk/tDYJ5K+AtvO
KoGYlkplvAXv1URN51GGq/Bp7fOVL5Zv7qbJ92CmqUEvqGuutB5qflchayFcS1xrQ7ukEfA58C4p
rmiwROAWrUD2K5pZZWO9AYQQYSsXXoZMYhakTINMp1SUbIfZO0NB1WHRn7SbhLh4GG5frdekUIfy
UC1Sh5oedymayvZpbe9wZDK74ZG/6kVG1HpFYtzrfZiG6+zgPtID979jtfkx3E6FCzGtDzksW9Q0
sqekIQIsrsi/n2SU1Rm4+nboWcYNykzisI+mP0T6MGvkTJs0wQL3XFE8KJ9QAL7ar/5SMKdURH2E
MXr8f/TzPGIYGGvkxbcMNw/04BnxkEpFfBQ6VHqFRM1cakbIhGJzgEoIrx8xB8Lz9uX0wEq0oJgK
/3CxUhiz0rRV8bLUYtUtgNgHCIa2qIz/lCQquos97slEAHWjfTrPzTs3Qx5a8hDtt3OLVTsDC4UB
sGj7DwuU4dDI2IA6lSWo012vkEe3xy9BxnwQT1zDJkF5+yWmOnogEMQMBtDMuSUzFCriCz03DOkh
wr2KSd/AXycWUmdrXl9YrCHOS722bF+nPAhJ2cx/CYiw2E8BY+mcU9vk74El+iHTGeqPWjBpDyP3
n3uCVgvzIJLer6TfCahSkjPim3P0QtYMRKGqjbqgpQ62Ffpttow+dneG2Sh50NxvZSKH1OAPA78P
D894+1Cb2ZrhjXqgnMptUlEKSQVJ4aaDyRF9klbteaJztKngTszfccxZVnm2DgKkRxDBOcnWDHyE
MCPH8UawA+hJt+rMXtITeybudmc05i9gbbfC/nWrVCDjEPup/QVjpwYLFYS3X8iOKRBhW6YkPa9N
vwosUUtEUc4oB9oRxe5RPNATWx/U2PSg2/yIruMIbvFVRImzuUTttcyI04D6lbgsAdgNoDWPOuMR
LP1S2HttNsP24Fk3PuIlgz8dNJU/SLcnGvazhgbyWWMMuIiF75TlK34oGJmBs75ax0IW9exvWXN8
Xlg2q+a9WVK1a09s+9FKMffJUrWFYdUS1/D7qek3klV8f0W5oVRjsYb4b+jGiBb8hD0RLaEMQciQ
QmyHYnPk39rbuLlyhMDEp6SIRkZvBbUisJCM5ZAjhcYapzgnHInw+NJV0aJc9TMIVRNv7aBDhi44
AwkIGRdM3+OGnRnVv71FzjMS2qTpaHtlZWjDkST12jgyYwx+lA5x2/R6c3XWxxrDTh2LaqPtBKHk
8LcDSOxwgF25RcMk2quXBaeYFwUTSPTLR+y4leQCTfxPu2Oxd18+PNoTojvEonPFCnN8ssYYFMvu
hKGGuC9ICsQTf/AvR7hS6kR8HqQljZTxqtwiIByDzs16t67yy63pNYij5goczLovvg7STTeNFdq4
ZBcVSLmDf02xXDrdZ85zGUv4hnWWnBOkFd4Y+euv3vgmcmutGwJtG2SLYprDbIOHLDVX/FJwxHiC
oDol9g1YO79ZrrbVF7o6vgChGHFOMa3TVRQOvVKuexslhNtkQK/X2dNI5P/ump+CDaZQPOEoKF68
FbsCRlxd6Uw1+TSPWAsQLP8KKskk4cZPcoASooG3tGnZUcOQnXUmVx7MH+fbPL4JBgcJOSPVCZ0J
CzxKzfRASbQS1MxEm55AY+ZF0I7TyBX577QjZDKXTXb2Gbqhm++pOXeWxUBSxYBBKg4IXNwkNabZ
8+D1fPN6oEyJoy/I1f/1CgRQBPgxM8BZ742Wz9XB7Twh9SvZx4uhu54pFfJEdSpM7lXWQIZYFsw6
gIRBsLl+HCI76xP1soshJQLGQbZXvpgqB9fZy3xEow/o1987wKt/jO5keogMBNZcOWgosd4tI1+V
eQmO9urRQABJE2gxfrlAT6bqQW4sCW6KGX70hF4PpC8dtGRzcis+va7b0UbjWg2Q3Ts63YYkCZoT
MbX98BT6sUFVyekgNSKm8dHR/cE2KJEKGcnlvIkgZn0u5ZjQAIcEVDszgdoKqM5bwxlqjeM6679e
6MyvevNQtE74jrKbimyMmkDhntdp/YtuYdMSAeu88bzN9AbMZ1WQ4JiiKvFMh07SnFSXdWLpZOFs
2a7n37Z2vZgQbYliXBFPx/mPOrIMh/giU3jqkOBLsXLqaxK4hylKJwQKXQmi36Ne8cL8fWFfVa4X
1rb09Df+uXjme+WD2Na2nPtUroVGarmpCmRqyw+PPMoQOnCwAowN0Xp14Zu5McizH8kJVZBAlcIN
m30o1rPr0ZgeJzslmEToGSEjHJdX1hHB/03Wo+HsNE1bs93ufjcDpQjeA56VBLZ0/1RQ3vd66Rr8
ZqdVHnRMCMyQ8OlRqAQFFlHdr632WK1g8Yq08gv/SIK/jCzBSaFc3FPfmhFazHVxTCZx+Ladbfph
6dLfAFduQj2RxZY0Foa+d7E6DmDdQLN7aBUfVBos4R3BupLInycho8lYGZN3dk5CJyi6VOXCDFG9
nvtn6KhH26kDb6taUk46YKAVSwZsXe9KauUVUGxinOGvqbb6D1MU7BL48Ymyxsxh9x9VXaWwzl2q
K8et8UZ0Ahf6bMI28fH4nNDn6KuxFao5l0PNt48Xjuvwe/v7by8FnlszrofPSWQrJ0XM2hmvINyW
+HxKyFlEi1EDjnr+wBp67EfSGKniqxlwscZlUi4yvYeP4VZt238RO+bW9uJkXPCslK4SGTfA14NQ
JmCdgaoFWbQehwS4SJrt/6C+M8/6H4SwegOs8pya0XmIfwbgQrzqBZPrZuw074uLo0wHenkdM0SN
AszP/4fZM2PF6s0H1CR93DEfeAu1JwRwvx3ZWMU5KdTlnSmpDrMyKAnMt7NA/QGlr0EvlZGlpUw0
naiiIPHKrcy1jXnmHbrY5QZi06w44QQhJMJUsr+clepSH7JArw1EMIIHwFr37C5oqFwXS22lFu2f
cCMiKitf91TVVGRwh+AUngG89Haxixb1mH78m5GCRLFsA+Pm9OMebbcPD9j2KTIv0L4Y6tX6RTCM
iqRXfATuapDrcssPoNTM0s0L2qIpBP5qCJLgPDflcPOllRgYcKziV5bgd09HouRamg9MfJ8oCEtF
QOSSdfcpdy0aaEhrwC0MA2DUQ0xlboDKCs/Sd1GKAKsdR+d+99ve/YW+Z90jfAWs5jkqS4+S9ARb
Yn/69yzskDYXCaHKTj3851VElAgZL5n1nzyaHef+G0lAZgfljYNTx4IhIL/oTsPYjwoAFNVTPXeD
Q+wm5dimB9qxbz9OIJxl/pNOftZifiXtluxUTEyCfytcSfNdmlXRCSf/OpLO88vBFs2ZE/oDwEob
CTia+6X/wYvZm6qdFgLJzZzMA8yZSofvDjrQMqfX8PbO2Kfu52s3v68BuNgteypURVIPr8zBlqgW
A6C5zRy0XR74bYtKSn/SVhhWhLAGI5m8bk13ef1EG1EF6Iy5JfLr6BxT5zGku4hIsdSp6l6s56zs
T1gpqLTlj6mxsBASPdfirnlAWiqsbHLBP8UZ4LRP8d5DT3pb5xEuJusGiRMwiZz2XdcacgrrHcIY
WZ37PvkYgwKxIX4yyXogvAD7+J3Uk7C/5kJgj/dAHH0HZNrAc+Ftw0g15Rz7ePANSI/X6bxt5lvJ
qhMwSM47Xq25q3pNil0kmKufJjpLHJHq7d7rILgkiYXbcw1ercP3fEV7MUuImlZWdTTECQVfrPy3
zc0qVkW1uymj0EqhaJM1a5raM48TvpKf3JRDjnr98ehfVS2OBp1R15QzrUWFHKrHCHw8GGSGfPma
ekGgLpkcy/6cGw6miP2x6CBlzT/NUeU+xiInxhcoaXkEig5SHn1w7vxh8E6yb9EurY8+NO41+FAZ
w1MHDe6Ed7KsIN/rgpFytVipWGbh1wHHHThi8xnyblSYEwf3m9x/xNj/hnBV6TW2Yd7J/0+74d2K
ID6K+IkfYTlvKe3/l3J6pcSl9Fk93pXt2k8S1yRnQqaiVJdTAcuJetPr6VPb9Ef6MW3iphA8h+Gu
vGiHNuyQpAFssfiiGq10k8ZarrRj/T5RdJJy7fueR9L3TeTe1SYQiCiELWxhcjmNMsnKKPX1sKof
/ZpYHKrNevVlAFBtfD7BX/1HL4c+C4BGJHiBCrsO2ilrPqWY8uLDyj/W+/oAfZCaNoA4kp+34PC4
gnSNC7EzWGJa8dmL41g02dEANGH2QEC8/eXB1aq5um25LTzA8JlZsMeJvmDwchkGVPOE8LR8pI0n
2EkpCVZp124HJ7AO7mrOj8kRKT5hT4IWJq6Fg6gVnXPC4K4j+NzrIXT3YaN1s9x5DZ1AAjkwvJz3
Bcjoit1tYbiqKS5V/+TUve+ziU8Dl+ymdevJ+/7sJ2O6zODEnpqRiUG81JlWlg5FiXr/p2zZINQH
vQtOQuTHh5oDqnRER/WLWaph4a6lVioxamzz0BhKPt5Y+3QKOMX9AWJCTmm0+FypJkfpNGvS8lld
DBJa2/NEBdy6Mt5U9cAkrvu75o+JOSJGQwa3F/GZbm/FJdg3NYnOzKSuxkiA+VFRfLBQwmcJE+MO
zJRpeb6qP+IgyMIP3Wxx9KPq2PfWb40eOHIVR8Q3VWaiuR5wHqmuEAC4I22UsTx2k2O4P6oLJbYj
ntaLKeE1jMFnS5pPtuL+HhiuVakPwi2pbFRN+QUHXxW9qmQzutTZgyz3W7mPKL40f0q5uQfFZhPV
Ze7JDadknuWmhSRgfrjNe6KaWYZQzyhQTVR4DC+SN7ZjsPaJXCNC391xt0ADRGgcI8XKdh30xuya
wgJnunWhYeFcf7USApGdrVqoSvr5q/JV/D7Z/N9L0P1LtSzphJBrsmLvGIv5oC5QHlSDQJLxH09q
rGygy+Ss4C8F8sgSt80HvqQG+NrsqxOTg9IQR00EfiFnQeR7WXATuVHU0KkQ1QUSpL6fbCZ8ywhe
qzF04zoF+QMC/R7vuOBWvfdKq0t8JmYE9oD7sc+iOeEccOhPuGXWVB07FRNHg51+l0Jv7R4eRoo8
R+lrQ/itEYxTgnS8zoflP1mV2GtSFUfIDHLxFFYfe254naetAl+wnHfNyVLG9nl8Kw2DhJomP20Z
czMrvjcTBQFc/hN1RgKvR/tCDVVkItDNvekMSEi+YAJ8iiHRKxMbcKeZr+a2k9ldepstk/RYUTyk
645wvD5tZiT+MJmSln/0svlLKQ0JmjDrMx8cHYHq4As1WDpAWhQbvLoJs3oCcDkTSSyt7USCiHU/
N6ZfcX4dqRJ5G2PVgOE2IEfWQY8FQ1qwBfv+dUUyH3N1KDQxsKNQSbsM1REVwLexqWcFmz0Gwq5P
7cg9ukZMjh0JHINU/ERTk2Z8coM4oUWJt6IT5X/CtzcNJcAQwFYY8Zo39pOvWItoI7epkHeEVTlp
3jMBHvPXS11pksQa86HNk3NCHG3FqLKNPuQk+KVAhn/oYr0dmwVMLVypUuWVfuGMehQU2T7Vv3wq
83LptX8x7sD3ftqAkmtPKYDFiUm+GAK4++8NPFe1tUtQdrK8ZsJb2zXa+qx3Ydp2HzhPJMUl8vE0
0Zk+M0lYQabEfo26QJPPT1jn1e4tSor7QCs5GuhSAMJxeFI5aUp7OeJlS1mpb4E89Pralm57WI7N
sScSosQKMUnfNL+QeipTSzu2X1GJ7UDvTGa+6a4VKEpdX1D0embCV1N36TYv19uDbApkjGA3mp9i
BcLhTvLZ6Oe0xiyx+OS76xw5/7H8f8KhjRQ5CWZ/WzVstFrC78VGS79PUGCQQqfIxZJOsBI0V0N6
hJkK+GhEwI1Axfp6SGfDCcPjMAf0CoRY9lh2pNDDugxaIzDkUfIeDUAHM/DGIpCS7/BOiFTzqRpJ
0NhIxAyPqxwEGnNqlPK/vMWpZ3D2TyPnulEn3jBCygH1oD8zqql99yItne4pW8+QOd7pmAEbx+Y4
7x7ukIbCCqjqVmW1u0Szl8+4VNU4damXbPS62rBf3bRcRTUK2P3nVU+x3Jcr20i7vK3KJv/kF5Yc
cBKKvf+KDgF+BtNl8k318Yh5jQ/Jh3Brv0LU+RIdSCZp/CvkbgklqS5ZslWM8+SrO9odfyflXUqr
hTsRpkDT67UtTScZfFzZu4vn/X3jdO0Xc/EZelKdvvDmTxrStwVvUKyP9REBsbHIzaTwZi+y+tPM
X2b4pvfx+Bh43e4FUkDAVPdipbUeMMnfsIaKJZNazlYm5JLNQ1hXZWZpBiY3VLXnOmZ2/pU8Pi/Y
i0StYiVcvJEpBGmpuJH7Jau62xQfEImmDnu1nNATDol8iRUbc/QoPhCbq3uhxDVC3r2vQlU0M+7V
Pn3PofZNsqLHL5JVhDOBF7LfQCu/PtyC9g/309p04OWvVIn26w8/k0o7FlxKLMMu1p2Vc+1Z9MkU
8BP7VWyK/lsdSRrKstESI93fWi2tCyfH90fLaXbZcqj2sYxx6B5px6xDldkerl1ql21GA0+nufG3
vWg9fay3LEYSGPNs+2fouogNQKIYjg6T56CLJ1PdVgbBHEcKwVhr73sjiCvr4cBNFaIPhdKUUEBK
QJFEtvSb0HEPhD69zlOGazJSGpmL/1oSKqsCbXDcbIj/m83OwKG16vTdwZo+weWH3vLClItryg3H
I0ctSfnqHlMozgFbsyF49Yi998R5QRakrBHWFdyDbJtKdqLu27KCdYMAsS4w21s7H7pbJePKPIuX
da6JpeOUHGZXpSJ7TxuSrWQDunq9EvXyrA6S8Xb6NnEVOh9Ryg/LTI//zwUBhko+qsHG86mysb2r
IQ/6z1I3htII/r1N0TR9fyGCo2+MsT3fCZXJ3Mq5bF86AxyiilM+NxhzDMZzaNiKDHe1CLCF/EI/
LwV6DM9thuTGo9P+rbnDs0v4ofdYby0/XAX3S40fUYiLXnscaIsXVKDP0KGe+z4YJOuMcYZO733V
I1YN258ImGrKWdhj9jxGu43SZRllVFfRxOsFbArT1+wyshdT+xCGB9vy9/mZ7Sja7IJu+O1sF+8b
lhcZ4iY/DPJlvDJI79jqgEb4LXNwI3tm4601YVsRi9nfMO5DGEIe4LfGjUpYTX9WAFUt7+7G3++T
+8HrXf7WJC3SeIEQJ3qKS/E+Z9kQxQt/0BodYF8Kf6+t1kfDW+LmFp+7OYH75kIy8DSaUqxNofrK
OTvPeWo+70mOxXq5vifG2oa95zgfaQN720FJWvnQ9uQGm70aHlGl5jSQ5yEUDSV1G4yUWSqQbodc
IcYNX8yhdVIxfUq44I5sBOiALSV1mRCXc4GafmyKYmFWMDHi5NVLcAiKa1+HeEPUWNsHa84sosKb
6KgNmUmJ/K9h20S1P1ty5Fs2TV15i4CjxaSZznmr9f/kAE1Okg1/e3W6/p/Qsy8PrUqCNlu7uNl2
hyMVru3roARDpD+XBQwF8SiAd8oePQPboTizqa2btsXoosMVbPrklpYpxkBegM9rOHYr3m3dEHpi
7htLi170ds9rhM1sE2g4kEToBbMedoKLrnjiOgCcIuj5kOFPPrhABnaTL3DAw+NTZt79QDEOCvBg
sa3ErSW6HB4VIRqq2zPjatgRlkLF3nvmRqzJn8NWK1kIHLJMU8E4OVRz+xp+NzQO5n5F4FmmCpAC
xE8IkyuUUPnfUtnfqexBeY03AQvHHXXvpi408xh//NxoI8mDxWimBbRTXhWYYxoJE9TKf33ec0NT
MZstvYcMVLBgR8Nc+Qi0B4FGn+6DlPr8PjDFowMWu0uH/qD3NDZkJGqNGNNgsjGm4psV2Dk/+rq9
wuOP8tI6CLYTaKTBddvnnu7k8XYputA6NYnqp5+TF3zlWGrrih+2wUYOHeWhq0Hk2fJAFeW/7mPK
+//iIwvwd/8Ux6yRq6RxKQWpsN3/FstxfvZE7FjNEKnCEDo018VbSksu3S3q0zOoWsCzmnpbUhEd
s5/Eot7XGlPeiZgIHL9lmer6oEuJGI7nf+aP/A3nFHUSPxEx5COY9Qik+PMqOpZDqIH7j42xewbs
Jq2rtb+35lxCL19zBxYxnHU87F5T9pnGAeQhSbO88Gix1cwMj55vTFY1njcMgOiEyX2eTt1UbAR2
ZhRz4MSnux7rRHLLbmZ+TDt2Gr+c2WJZMrUCZw31fEv6AyR2upHJ+e343nzBthGsGl3w1yzQhx6u
XJCbsRGDjfoouRyRnPCRJGUqThwQl4+Cb+6AYE0pg8wKT12AoNShejv9xL0L/3T7V0lSXwbj7lyO
PYhyxBydIsg83pEaKHZuwkFBGgiJBPQmSx/EX4pikR1fgBpQgyHcc901cbdADeohq2p6xd6gsPHt
JnH012SDq2OhQvWwDTEQwcqual19EqwgFreEKFKeceaOE4Zr0qo55YpvLWnecIpcz0G9mQPmYnVt
UoPETuTiVX4CnjtDpie7t1Yezu9Z+GL7jfpkix0Srrmm/yDtij6RZCjACVo+qRxzQscM3BZzHiMw
z1gWDIQLnog5P5IHpliU5bmGIy6Kwt8FxRr38tPdI+ExE3VrzWmTdnT59O7/ZGvmIuWRny/wqDff
uEo876F+oNSY57UJfLqHZ1nalbrPNW1oakjoFKo5tghgov+XkCsJt5yEHWq9m7+uM/I04c8Y01f0
3ngNtYl0JTbgGiK70SGifPEyQAUmeLHRzfPJDM6PnkT+jWPc/qdGJM4V3AqyIKkV18gwbQuu7K9S
P7xynEyuExy4gBR+YRvj19tr9bIlifXvQRyu2WFG9tV/RWR8xS+fYLhonl0SPs6vqfIvx5v52DRT
a6jWfQqqMT5bqUXFwzuqw0SEpYYrojzzIkpc5DlVx2VGmYnZvle+/VkHZE8LO012+0EMLARFRy/w
DsUmBrXVO89K5PqroKYvSPDG6YLE2xR+sxxG5nW30HMDQf8NSZ2G8c3RJ8o7x/lQBq1sTK+Hxsvx
D4HhSKOnx7ACPNQ4SvwW6X0pDGlMiRUTdAnfjoaUh0PivHD03AmRmtG9RkTkDwFi0RIR40oH3q91
V55lsGayDfXjAvCVZvagM/U+swLisle7SFRgyd5TkUvALLnljJJWYNorN/hJ/FfIxyc9IT27v5xC
MGciILcaU5OXtxek8//9rORcjAOje81l6ps3G2LJZzQhcPWPldVVZ+8Ia3rzCkWlTZJo9wNCmBUr
vgkLIxt8ewb1U3IZnmPDqvjoBIYLdLkKNYSqj4v6BvFEdkMbbsZg9uX8o6VsDiUUKraqkWA6nQld
JvclgBXmtSASyf5SE3rhQbnD8vpDHuertzwkYUQzWVVQyeSqbyQafMrnkpfFwphTtI6TvN7dLkMJ
ka3yj1r49iWtPyNnHlay3Bbq9cri0N0KQFjxamYFSnmcGyL8JOUZqh4FEUS0TEOVDF+RdUKmKmNR
LRtEvL+5BTH5aQsNwJfKO2KPUsuWNgqgrvrXpC0B5o9UaGNA8IVD/16BVlv2QfqPqYhasQLDd29A
D41m4NjVtH09kRCR5p2toubhHrIEOdWpltcPbVaI/8XXrMq5OESrhF91cmvb7YoJuw2bMqV1LClg
5WDYEN1D0BL5qxsUvixPd6eLAKtfQG4xjqOnY12q8KbkrD16fxge3as1hvMnsN0PkY/ZNlM0cOhg
9OjjG0snIet+ZQv9ZTGeIfRB87wWJ8Rd0ye7BSGcDyYe1aYq6bvCAJX39g6G9tlMm6dmIp2MY6pF
mGYlBsQ8TmDNwcu+jTbwzoAwFWeO3XDyMVPjtExZ8d+sGuQu7Gqxff8GQWnT8Mn1vvVbIlWamR1W
nvWHvWnMJiv3l0j4LdovjmcVQFbPMQ9uE33Ks0vswCib5LUvta5k9Ml0c/jUSmSbRpKxaSIa1QI2
/uu2qWvFbQhrnXAF7n2n+KeVrpB8G1dXfpzkKWPZHzWp6suiLOQ4atzk7F+NYp0wzDqdB3Wx/uWo
eHZsTctfWwHpVTEkHU9Yex3QAuFd2GX95iVElHgw/7zSe0s9xJTten291MO3HCim/RQbNxKad7Am
HbS/OE+dmiURIfdXRaqlBGiYFg4uWHVp0eYWM1MonGPpQFIJEpZlyijmgxs7x75JZwS4KGEIJ25i
mlYxSon2Qm7ZaNkEPJPA4SU/e9I8fVyU23ByCNYrxalcme+rFOPuzlFMD34YkcsxywsDYfyptTaw
Ii2u4lXuVldNPd8NYyYoxwxUGC9MGd8gaIpFjtgrffFCDT6lC3z3hDZ1IfIOiLwwljrW9IxsjMo8
9JKjqJu2h2sJVeiXCdFH8ElGBfZXVl2SG+yV3eVUUrao5els2wa1K5iTkhVi3sGWK1huQiVITGR+
Ea0tacwaPi+k4bTW/7A68E0RBvW/qqImn5OeB+sHfSzHyQQi+Hm5FXpCD7LFiIGtmh3uphc7PIlq
sc31BWEE/DGxU2us7cd0hMBcHjMKj8/6lFJ9fCUrJsDHrvSJv7cyekc5P9MnxIixSI2b2pLoJXWN
MbNnukk+gqsYlWf6+VYFeZrm32MQFjxx0/6jtuah0cRTPmy8oeHOAtjFOX4SIPvLOREbVq9REURr
z2tP2qCUUGukFvsrgUpJQE6kq3mfJZxyoTUJG8LUtuZAovtKkKfZqVrlXN2TCk6jpaAJBzO3HWNX
Z1hogUYVdjHOP/vtEkG4le3ZoF5dou9XS+Uy2H8HuR1T/p9kA4CnT+7YOmZrxj9IEj6nFg3adnjx
ClChkRys3FkB4LSCXySb7O5Xvwh+o9ORpYLn9/UDy+ZM04kiddRL9qj94GghhRWV792vmQVUFa/B
Qi20ufHJArDKO9ZmQv0nYnOmeGVxrSt3eDZXC4CJuoZFeOhG2hMYyRk63mvRRVbyvp7kRZ2H6GUx
Jdr7UaA34bQbTCpnYIlCAbn5xtFOWzC5THLagnMy330K44Kq0IroMDbRvPLIg9HJfKSipI7S9kT4
42kXEf1koFG+p9sru3J41ig30dhmvtecdQuVEGkvcq8GdluKK/5uVqxyINg/pLvNV+2Tj11W6lfQ
LEg0ds6a2zayTJLTtPQo5UCApZqohBYDR4OKv7tV6EuZw6YhMTsTG9auhsma+Rvm3GfpNsw3SJpQ
6t+25HYB2y78PANb8nVtbNnpjKa3ZpWUnHGEjprcQhq3gsz59llt1rUI77eQMlT0X7KTq5y3IUxQ
i54XICNIWs+e2FaiyNfMZMNn/979kaC8f0/iwAs/ITmCPOmg8cD1nXu6/4xGvur77J08VmM/yxHP
6gsG/0jNb9dzJ7reBJZzHPurZaKtGfnPCm6GIXiT6xmWGqc8MD6HtvwLfGfV3/431/GRL9PnhdRY
dpqKRJLvcH4HHNXuTDCCCEc4Ic8TSXI5XWSAsFf97Sm99k4F9d5g1IMxFJVLVDEbBhhhjD1BWgMB
bEDob7iy6FCiTfTvAIjzRgI6S6Bn4YewQiqbFvABKq1Nkqt4/+z6vaDZRfD7lOH3F6rod39vFznD
o37bELMV6RSnDI280NH7+XKK5KpFms7j5Dl1Vc14SbssMH/sdOHOuOUKtg4S6gU5UewKK4TI9KP0
tADCztJ8UqCpG2FyEtcIwA8ASpQV/40sLIshRyuLwL7sv3pDFsNGI1VH8bIY1PAHbBve8oZZ7JhJ
9D2ng/VXMf6TDnkCywVmpkWm7M46HZfRAMjQ+QYbGCEPyBQNsam3zraiRkm61dwegfY3GVu6CS6S
tJHAcysW93CfwQDefon+C1ZENrU3mykwmJmCzLtvOc7+MxVxy5lruN2vJSsJalZUoFsHjr15X2aV
cmGCuLuedsCD+F7x7zutaCTP9++tsYpZiLfCNrhIHzwTxiFyw/cGmkxBj8LcmpIRDsXucatC1Kpm
noXsEriCgO5i47V/AGJBaVl+VdH+1sYbpm8NC5l5QejCVaE0EjElambLhcjVn03WkvBh4dL3BREx
OfGW71NWMNvBS/Npvuw5KS//zKgx0qTrr+zquXjdjkJeKZDkjWcX2wxPlIDt2LAqlUxecAyacZqX
fdH8ou2dkAX8fFlB0L0Sr6i8p2fRkdFCKu72wAY0ej4ZgNrlf8cTIj7vR1BCDCOdi9T3lLyfWD7A
Px0lowR0989Dka/rGpc6otCCEEwxmvKsh8kCfmLvmOKpAtUoWXw3V8KcGrOQwXEDIdkiVvzI7Kva
rhfgc18E+M/x9sBVWGaQ/3jjR/AyL5Q6zweS/PH5DxIO+gp3Ao0uxzXLFs/Gry6m2K3oYZ5dQRMu
pjwE0yLIOaexboCLQFIDHfb+Ga9ckQJ9g/v4oqi5TP37NmjH26stbZmZvQE1LFoLinFidNj2xVdY
uDRsOgfbSwyueDcerLZ2k6OvWY+RgQ1++v4+rgons8cbTVFmOuhVlQeQa6k+JS13HFIm8vZNDCRC
fgl1duH0S0oDzAyN44hBWT6j9D97Ur+uN3u8abg2qOYPmQezG004PqagMhEQv+tTM/N8a3H29C1n
+gME+MT4A+JnobHiDBpIQp0HsZQkM1b/n4W3KrFh7+Nfi2mGFEzusd6Dh1ZCzr5ri/MIMQZVJo3P
zU4qTDvgpswy+ZNuCHbCBNXvIpSnSZFTsi0H9E7XynF4cRdjb+xHnXtxl0PHVemhsRL9Tb7fpu3V
PaHtRxVX8drJMP+ZYKRaMArcS9+914dETYOzQp94N2R+kXXgSQsT2480CUfclXEN9fc1L4YkCa6/
rZHOa9jL6J8O3neDaW0BS6ZGpp3+OWCJz2lJ9bGpNikTGz/049X2CEneyMSMPwHCofgmqC+yxp8b
9Mp+E0KJKrVeTa3OThgxw6WldvOyHyxt0hvKMjJ0QOgmvtWywAjc4KCWmyc/aa//9k2Ao+5QTVxe
hEjt/jQN+4N87/CMMF9fOxUy8N98Snq9gzeE/XQsDcHaJ5r4G1dEwmzN6iMYAt0W+i3+fbekY/Qa
J0zbhR+nTPhdjX3w41rqv8yTSJsw6+jFYJJii8RUsjfWAdYO//Sjufl++qM8ks4ILNWkMEobq0z6
FWM4qW0FZ8OQm90ey7O7bsuOxgcNzO6+0GQu1XEr5wwFgSCHnMbUjlrl40J4U3mhyOUU8FHmJLZa
f+jV+aPx5tyBrrSzQvEvpRAR7CGijnU2H7I+5UPXqZa5PUCyiHJYCgOiJBqGJJ0/HYJWDzm6kfhx
G5iPCHt7chalIp5dYRjHEX9gLWKMcDhrbiDkyp9u+AnEPRfUyRRKz1jew12PeWiITdf4p9qYg0Lt
e0b5+5t+lDJr/5qshCK1h0QnXREYHQN6YeUQol56SCN19ESU7mWfvKD0PEd+YkvFOExGIH9xOd/i
nuq4CqzmBnpG5ZkL0yPI0veTBut3WHOThy56q0Vy0ht/PbVXzgiNs9GgSlPPQSLeWnhi3pz91G+5
f/MqfnT/me5fcP5vabxRnTU0hXRs4XAlmvg8uR2TdZZQnLHgQRguojo334u1myPSLXbA+Aizsp7I
z0+UZFoNfZBCCLGQhJSl+qE8AVq5xb8ry/NM54iXWlLVEVKasOWB/7ytR/boBL+dv87V6BO8TeoH
fCvP6WsLrFX0HNTynr84+KkUkogB559wQo6kk5IPXWZoeFDxGMSfrT+PcgkxGGyH02azrMENDU0a
U4V3+yoSRfFOTR/e8s4Tqhvzjz4XC06WkpDq14wIRD+rG8BstdUE3nI7d3Z4zTgpm5MYJupAdNNl
YQ5qVZnidzWRYRWFqB/cHj3bTJ4UurOdSSJs/j7lZ5GexwVJqaL5tO5wjcyRxh5WbmhZYi1+gh7g
o8LlFLjowaLYkjmEWZM0Cx9RKfWEUQ9GW3jSSRxN7u7ahAqazxbwOnxz7NVx94Yu2yDq0BP+Ie+Z
70lPLaX5d4Kphe6Bd4/vDo8O29KsNySvMMWlze+uQRhsQNtaula9nxrJqDw5kbPdi8toN7OwN+Ss
4oPklpn3ddNeZhrcXeOcYSDp7QlJdZ+1J5y4ZLgt0fyTzHxw1rvCNRQQVmjBaaJMvCen3n8QzJ5v
MvUy+yotxOcBeOouIN1g/P7jH6u7abe1vj7Ofpt+tP+NLXjFYPezoTZc+tB5+3eQBu8=
`protect end_protected
