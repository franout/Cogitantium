// Register NVDLA_CFGROM_CFGROM_HW_VERSION_0
#define NVDLA_CFGROM_CFGROM_HW_VERSION_0					32'h0
#define NVDLA_CFGROM_CFGROM_HW_VERSION_0_HW_VERSION_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_HW_VERSION_0_HW_VERSION_SIZE				32


// Register NVDLA_CFGROM_CFGROM_GLB_DESC_0
#define NVDLA_CFGROM_CFGROM_GLB_DESC_0					32'h4
#define NVDLA_CFGROM_CFGROM_GLB_DESC_0_GLB_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_GLB_DESC_0_GLB_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_DESC_0
#define NVDLA_CFGROM_CFGROM_CIF_DESC_0					32'h8
#define NVDLA_CFGROM_CFGROM_CIF_DESC_0_CIF_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_DESC_0_CIF_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0					32'hc
#define NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0_CIF_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0_CIF_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0					32'h10
#define NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0_CIF_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0_CIF_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0					32'h14
#define NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0_CIF_BASE_WIDTH_RANGE			7:0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0_CIF_BASE_WIDTH_SIZE				8


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0					32'h18
#define NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0_CIF_BASE_LATENCY_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0_CIF_BASE_LATENCY_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0					32'h1c
#define NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0_BASE_BURST_LENGTH_MAX_RANGE			31:5
#define NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0_BASE_BURST_LENGTH_MAX_SIZE				27


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0					32'h20
#define NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0_CIF_BASE_MEM_ADDR_WIDTH_RANGE			31:5
#define NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0_CIF_BASE_MEM_ADDR_WIDTH_SIZE				27


// Register NVDLA_CFGROM_CFGROM_CDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_CDMA_DESC_0					32'h24
#define NVDLA_CFGROM_CFGROM_CDMA_DESC_0_CDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_DESC_0_CDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0					32'h28
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0_CDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0_CDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0					32'h2c
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0_CDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0_CDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0					32'h30
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0_CDMA_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0_CDMA_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0					32'h34
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0_CDMA_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0_CDMA_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0					32'h38
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0_CDMA_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0_CDMA_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0					32'h3c
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0_CDMA_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0_CDMA_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0					32'h40
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0_CDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0_CDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0					32'h44
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0_CDMA_BASE_CBUF_BANK_NUM_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0_CDMA_BASE_CBUF_BANK_NUM_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0					32'h48
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0_CDMA_BASE_CBUF_BANK_WIDTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0_CDMA_BASE_CBUF_BANK_WIDTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0					32'h4c
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0_CDMA_BASE_CBUF_BANK_DEPTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0_CDMA_BASE_CBUF_BANK_DEPTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0					32'h50
#define NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0_CDMA_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0_CDMA_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0					32'h54
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0_CDMA_IMAGE_IN_FORMATS_PACKED_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0_CDMA_IMAGE_IN_FORMATS_PACKED_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0					32'h58
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0_CDMA_IMAGE_IN_FORMATS_SEMI_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0_CDMA_IMAGE_IN_FORMATS_SEMI_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_DESC_0
#define NVDLA_CFGROM_CFGROM_CBUF_DESC_0					32'h5c
#define NVDLA_CFGROM_CFGROM_CBUF_DESC_0_CBUF_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_DESC_0_CBUF_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0					32'h60
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0_CBUF_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0_CBUF_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0					32'h64
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0_CBUF_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0_CBUF_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0					32'h68
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0_CBUF_BASE_CBUF_BANK_NUM_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0_CBUF_BASE_CBUF_BANK_NUM_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0					32'h6c
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0_CBUF_BASE_CBUF_BANK_WIDTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0_CBUF_BASE_CBUF_BANK_WIDTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0					32'h70
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0_CBUF_BASE_CBUF_BANK_DEPTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0_CBUF_BASE_CBUF_BANK_DEPTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0					32'h74
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0_CBUF_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0_CBUF_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_DESC_0
#define NVDLA_CFGROM_CFGROM_CSC_DESC_0					32'h78
#define NVDLA_CFGROM_CFGROM_CSC_DESC_0_CSC_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_DESC_0_CSC_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0					32'h7c
#define NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0_CSC_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0_CSC_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0					32'h80
#define NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0_CSC_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0_CSC_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0					32'h84
#define NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0_CSC_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0_CSC_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0					32'h88
#define NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0_CSC_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0_CSC_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0					32'h8c
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0_CSC_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0_CSC_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0					32'h90
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0_CSC_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0_CSC_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0					32'h94
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0_CSC_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0_CSC_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0					32'h98
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0_CSC_BASE_CBUF_BANK_NUM_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0_CSC_BASE_CBUF_BANK_NUM_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0					32'h9c
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0_CSC_BASE_CBUF_BANK_WIDTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0_CSC_BASE_CBUF_BANK_WIDTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0					32'ha0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0_CSC_BASE_CBUF_BANK_DEPTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0_CSC_BASE_CBUF_BANK_DEPTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0					32'ha4
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0_CSC_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0_CSC_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0					32'ha8
#define NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0_CSC_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0_CSC_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0					32'hac
#define NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0_CMAC_A_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0_CMAC_A_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0					32'hb0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0_CMAC_A_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0_CMAC_A_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0					32'hb4
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0_CMAC_A_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0_CMAC_A_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0					32'hb8
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0_CMAC_A_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0_CMAC_A_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0					32'hbc
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0_CMAC_A_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0_CMAC_A_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0					32'hc0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0_CMAC_A_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0_CMAC_A_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0					32'hc4
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0_CMAC_A_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0_CMAC_A_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0					32'hc8
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0_CMAC_A_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0_CMAC_A_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0					32'hcc
#define NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0_CMAC_B_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0_CMAC_B_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0					32'hd0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0_CMAC_B_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0_CMAC_B_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0					32'hd4
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0_CMAC_B_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0_CMAC_B_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0					32'hd8
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0_CMAC_B_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0_CMAC_B_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0					32'hdc
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0_CMAC_B_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0_CMAC_B_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0					32'he0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0_CMAC_B_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0_CMAC_B_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0					32'he4
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0_CMAC_B_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0_CMAC_B_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0					32'he8
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0_CMAC_B_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0_CMAC_B_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_DESC_0
#define NVDLA_CFGROM_CFGROM_CACC_DESC_0					32'hec
#define NVDLA_CFGROM_CFGROM_CACC_DESC_0_CACC_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_DESC_0_CACC_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0					32'hf0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0_CACC_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0_CACC_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0					32'hf4
#define NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0_CACC_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0_CACC_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0					32'hf8
#define NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0_CACC_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0_CACC_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0					32'hfc
#define NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0_CACC_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0_CACC_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0					32'h100
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0_CACC_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0_CACC_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0					32'h104
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0_CACC_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0_CACC_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0					32'h108
#define NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0_CACC_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0_CACC_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0					32'h10c
#define NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0_CACC_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0_CACC_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0					32'h110
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0_SDP_RDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0_SDP_RDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0					32'h114
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0_SDP_RDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0_SDP_RDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0					32'h118
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0_SDP_RDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0_SDP_RDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0					32'h11c
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0_SDP_RDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0_SDP_RDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0					32'h120
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0_SDP_RDMA_BASE_SDP_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0_SDP_RDMA_BASE_SDP_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_DESC_0
#define NVDLA_CFGROM_CFGROM_SDP_DESC_0					32'h124
#define NVDLA_CFGROM_CFGROM_SDP_DESC_0_SDP_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_DESC_0_SDP_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0					32'h128
#define NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0_SDP_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0_SDP_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0					32'h12c
#define NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0_SDP_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0_SDP_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0					32'h130
#define NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0_SDP_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0_SDP_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0					32'h134
#define NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0_SDP_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0_SDP_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0					32'h138
#define NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0_SDP_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0_SDP_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0					32'h13c
#define NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0_SDP_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0_SDP_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0					32'h140
#define NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0_SDP_BS_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0_SDP_BS_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0					32'h144
#define NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0_SDP_BN_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0_SDP_BN_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0					32'h148
#define NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0_SDP_EW_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0_SDP_EW_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0					32'h14c
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0_PDP_RDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0_PDP_RDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0					32'h150
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0_PDP_RDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0_PDP_RDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0					32'h154
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0_PDP_RDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0_PDP_RDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0					32'h158
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0_PDP_RDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0_PDP_RDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0					32'h15c
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0_PDP_RDMA_BASE_PDP_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0_PDP_RDMA_BASE_PDP_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_DESC_0
#define NVDLA_CFGROM_CFGROM_PDP_DESC_0					32'h160
#define NVDLA_CFGROM_CFGROM_PDP_DESC_0_PDP_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_DESC_0_PDP_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0					32'h164
#define NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0_PDP_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0_PDP_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0					32'h168
#define NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0_PDP_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0_PDP_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0					32'h16c
#define NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0_PDP_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0_PDP_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0					32'h170
#define NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0_PDP_BASE_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0_PDP_BASE_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0					32'h174
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0_CDP_RDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0_CDP_RDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0					32'h178
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0_CDP_RDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0_CDP_RDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0					32'h17c
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0_CDP_RDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0_CDP_RDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0					32'h180
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0_CDP_RDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0_CDP_RDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0					32'h184
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0_CDP_RDMA_BASE_CDP_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0_CDP_RDMA_BASE_CDP_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_DESC_0
#define NVDLA_CFGROM_CFGROM_CDP_DESC_0					32'h188
#define NVDLA_CFGROM_CFGROM_CDP_DESC_0_CDP_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_DESC_0_CDP_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0					32'h18c
#define NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0_CDP_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0_CDP_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0					32'h190
#define NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0_CDP_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0_CDP_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0					32'h194
#define NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0_CDP_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0_CDP_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0					32'h198
#define NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0_CDP_BASE_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0_CDP_BASE_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_END_OF_LIST_0
#define NVDLA_CFGROM_CFGROM_END_OF_LIST_0					32'h19c
#define NVDLA_CFGROM_CFGROM_END_OF_LIST_0_END_OF_LIST_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_END_OF_LIST_0_END_OF_LIST_SIZE				32


// Register NVDLA_GLB_S_NVDLA_HW_VERSION_0
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0					32'h1000
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MAJOR_RANGE			7:0
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MAJOR_SIZE				8
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MINOR_RANGE			23:8
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MINOR_SIZE				16


// Register NVDLA_GLB_S_INTR_MASK_0
#define NVDLA_GLB_S_INTR_MASK_0					32'h1004
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK0_RANGE			0:0
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK1_RANGE			1:1
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK0_RANGE			2:2
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK1_RANGE			3:3
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK0_RANGE			4:4
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK1_RANGE			5:5
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK0_RANGE			6:6
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK1_RANGE			7:7
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK0_RANGE			8:8
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK1_RANGE			9:9
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK0_RANGE			16:16
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK1_RANGE			17:17
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK0_RANGE			18:18
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK1_RANGE			19:19
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK0_RANGE			20:20
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK1_RANGE			21:21
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK1_SIZE				1


// Register NVDLA_GLB_S_INTR_SET_0
#define NVDLA_GLB_S_INTR_SET_0					32'h1008
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET0_RANGE			0:0
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET1_RANGE			1:1
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET0_RANGE			2:2
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET1_RANGE			3:3
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET0_RANGE			4:4
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET1_RANGE			5:5
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET0_RANGE			6:6
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET1_RANGE			7:7
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET0_RANGE			8:8
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET1_RANGE			9:9
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET0_RANGE			16:16
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET1_RANGE			17:17
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET0_RANGE			18:18
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET1_RANGE			19:19
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET0_RANGE			20:20
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET1_RANGE			21:21
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET1_SIZE				1


// Register NVDLA_GLB_S_INTR_STATUS_0
#define NVDLA_GLB_S_INTR_STATUS_0					32'h100c
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS0_RANGE			0:0
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS1_RANGE			1:1
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS0_RANGE			2:2
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS1_RANGE			3:3
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS0_RANGE			4:4
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS1_RANGE			5:5
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS0_RANGE			6:6
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS1_RANGE			7:7
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS0_RANGE			8:8
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS1_RANGE			9:9
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS0_RANGE			16:16
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS1_RANGE			17:17
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS0_RANGE			18:18
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS1_RANGE			19:19
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS0_RANGE			20:20
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS1_RANGE			21:21
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS1_SIZE				1


// Register NVDLA_MCIF_CFG_RD_WEIGHT_0_0
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0					32'h2000
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_BDMA_RANGE			7:0
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_BDMA_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_SDP_RANGE			15:8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_SDP_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_PDP_RANGE			23:16
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_PDP_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_CDP_RANGE			31:24
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_CDP_SIZE				8


// Register NVDLA_MCIF_CFG_RD_WEIGHT_1_0
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0					32'h2004
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_B_RANGE			7:0
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_B_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_N_RANGE			15:8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_N_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_E_RANGE			23:16
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_E_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_CDMA_DAT_RANGE			31:24
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_CDMA_DAT_SIZE				8


// Register NVDLA_MCIF_CFG_RD_WEIGHT_2_0
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0					32'h2008
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_CDMA_WT_RANGE			7:0
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_CDMA_WT_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RBK_RANGE			15:8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RBK_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_1_RANGE			23:16
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_1_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_0_RANGE			31:24
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_0_SIZE				8


// Register NVDLA_MCIF_CFG_WR_WEIGHT_0_0
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0					32'h200c
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_BDMA_RANGE			7:0
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_BDMA_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_SDP_RANGE			15:8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_SDP_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_PDP_RANGE			23:16
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_PDP_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_CDP_RANGE			31:24
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_CDP_SIZE				8


// Register NVDLA_MCIF_CFG_WR_WEIGHT_1_0
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0					32'h2010
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RBK_RANGE			7:0
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RBK_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_2_RANGE			15:8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_2_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_1_RANGE			23:16
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_1_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_0_RANGE			31:24
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_0_SIZE				8


// Register NVDLA_MCIF_CFG_OUTSTANDING_CNT_0
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0					32'h2014
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_RD_OS_CNT_RANGE			7:0
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_RD_OS_CNT_SIZE				8
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_WR_OS_CNT_RANGE			15:8
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_WR_OS_CNT_SIZE				8


// Register NVDLA_MCIF_STATUS_0
#define NVDLA_MCIF_STATUS_0					32'h2018
#define NVDLA_MCIF_STATUS_0_IDLE_RANGE			8:8
#define NVDLA_MCIF_STATUS_0_IDLE_SIZE				1
#define NVDLA_MCIF_STATUS_0_IDLE_NO			1'h0
#define NVDLA_MCIF_STATUS_0_IDLE_YES			1'h1


// Register NVDLA_CDMA_S_STATUS_0
#define NVDLA_CDMA_S_STATUS_0					32'h3000
#define NVDLA_CDMA_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CDMA_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CDMA_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CDMA_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CDMA_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CDMA_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CDMA_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CDMA_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CDMA_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CDMA_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CDMA_S_POINTER_0
#define NVDLA_CDMA_S_POINTER_0					32'h3004
#define NVDLA_CDMA_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CDMA_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CDMA_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CDMA_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CDMA_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CDMA_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CDMA_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CDMA_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CDMA_S_ARBITER_0
#define NVDLA_CDMA_S_ARBITER_0					32'h3008
#define NVDLA_CDMA_S_ARBITER_0_ARB_WEIGHT_RANGE			3:0
#define NVDLA_CDMA_S_ARBITER_0_ARB_WEIGHT_SIZE				4
#define NVDLA_CDMA_S_ARBITER_0_ARB_WMB_RANGE			19:16
#define NVDLA_CDMA_S_ARBITER_0_ARB_WMB_SIZE				4


// Register NVDLA_CDMA_S_CBUF_FLUSH_STATUS_0
#define NVDLA_CDMA_S_CBUF_FLUSH_STATUS_0					32'h300c
#define NVDLA_CDMA_S_CBUF_FLUSH_STATUS_0_FLUSH_DONE_RANGE			0:0
#define NVDLA_CDMA_S_CBUF_FLUSH_STATUS_0_FLUSH_DONE_SIZE				1


// Register NVDLA_CDMA_D_OP_ENABLE_0
#define NVDLA_CDMA_D_OP_ENABLE_0					32'h3010
#define NVDLA_CDMA_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CDMA_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CDMA_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CDMA_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CDMA_D_MISC_CFG_0
#define NVDLA_CDMA_D_MISC_CFG_0					32'h3014
#define NVDLA_CDMA_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CDMA_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CDMA_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CDMA_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CDMA_D_MISC_CFG_0_IN_PRECISION_RANGE			9:8
#define NVDLA_CDMA_D_MISC_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_CDMA_D_MISC_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_CDMA_D_MISC_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_CDMA_D_MISC_CFG_0_IN_PRECISION_FP16			2'h2
#define NVDLA_CDMA_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CDMA_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CDMA_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CDMA_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CDMA_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_CDMA_D_MISC_CFG_0_DATA_REUSE_RANGE			16:16
#define NVDLA_CDMA_D_MISC_CFG_0_DATA_REUSE_SIZE				1
#define NVDLA_CDMA_D_MISC_CFG_0_DATA_REUSE_DISABLE			1'h0
#define NVDLA_CDMA_D_MISC_CFG_0_DATA_REUSE_ENABLE			1'h1
#define NVDLA_CDMA_D_MISC_CFG_0_WEIGHT_REUSE_RANGE			20:20
#define NVDLA_CDMA_D_MISC_CFG_0_WEIGHT_REUSE_SIZE				1
#define NVDLA_CDMA_D_MISC_CFG_0_WEIGHT_REUSE_DISABLE			1'h0
#define NVDLA_CDMA_D_MISC_CFG_0_WEIGHT_REUSE_ENABLE			1'h1
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_DATA_RLS_RANGE			24:24
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_DATA_RLS_SIZE				1
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_DATA_RLS_DISABLE			1'h0
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_DATA_RLS_ENABLE			1'h1
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_WEIGHT_RLS_RANGE			28:28
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_WEIGHT_RLS_SIZE				1
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_WEIGHT_RLS_DISABLE			1'h0
#define NVDLA_CDMA_D_MISC_CFG_0_SKIP_WEIGHT_RLS_ENABLE			1'h1


// Register NVDLA_CDMA_D_DATAIN_FORMAT_0
#define NVDLA_CDMA_D_DATAIN_FORMAT_0					32'h3018
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_DATAIN_FORMAT_RANGE			0:0
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_DATAIN_FORMAT_SIZE				1
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_DATAIN_FORMAT_FEATURE			1'h0
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_DATAIN_FORMAT_PIXEL			1'h1
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_RANGE			13:8
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_SIZE				6
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R8			6'h0
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R10			6'h1
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R12			6'h2
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R16			6'h3
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R16_I			6'h4
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R16_F			6'h5
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A16B16G16R16			6'h6
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_X16B16G16R16			6'h7
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A16B16G16R16_F			6'h8
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A16Y16U16V16			6'h9
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_V16U16Y16A16			6'ha
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A16Y16U16V16_F			6'hb
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A8B8G8R8			6'hc
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A8R8G8B8			6'hd
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_B8G8R8A8			6'he
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R8G8B8A8			6'hf
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_X8B8G8R8			6'h10
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_X8R8G8B8			6'h11
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_B8G8R8X8			6'h12
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R8G8B8X8			6'h13
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A2B10G10R10			6'h14
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A2R10G10B10			6'h15
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_B10G10R10A2			6'h16
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_R10G10B10A2			6'h17
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A2Y10U10V10			6'h18
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_V10U10Y10A2			6'h19
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_A8Y8U8V8			6'h1a
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_V8U8Y8A8			6'h1b
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y8___U8V8_N444			6'h1c
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y8___V8U8_N444			6'h1d
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y10___U10V10_N444			6'h1e
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y10___V10U10_N444			6'h1f
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y12___U12V12_N444			6'h20
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y12___V12U12_N444			6'h21
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y16___U16V16_N444			6'h22
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_FORMAT_T_Y16___V16U16_N444			6'h23
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_MAPPING_RANGE			16:16
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_MAPPING_SIZE				1
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_MAPPING_PITCH_LINEAR			1'h0
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_MAPPING_RESERVED_LINEAR			1'h1
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_SIGN_OVERRIDE_RANGE			20:20
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_SIGN_OVERRIDE_SIZE				1
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_SIGN_OVERRIDE_UNSIGNED_INT			1'h0
#define NVDLA_CDMA_D_DATAIN_FORMAT_0_PIXEL_SIGN_OVERRIDE_SIGNED_INT			1'h1


// Register NVDLA_CDMA_D_DATAIN_SIZE_0_0
#define NVDLA_CDMA_D_DATAIN_SIZE_0_0					32'h301c
#define NVDLA_CDMA_D_DATAIN_SIZE_0_0_DATAIN_WIDTH_RANGE			12:0
#define NVDLA_CDMA_D_DATAIN_SIZE_0_0_DATAIN_WIDTH_SIZE				13
#define NVDLA_CDMA_D_DATAIN_SIZE_0_0_DATAIN_HEIGHT_RANGE			28:16
#define NVDLA_CDMA_D_DATAIN_SIZE_0_0_DATAIN_HEIGHT_SIZE				13


// Register NVDLA_CDMA_D_DATAIN_SIZE_1_0
#define NVDLA_CDMA_D_DATAIN_SIZE_1_0					32'h3020
#define NVDLA_CDMA_D_DATAIN_SIZE_1_0_DATAIN_CHANNEL_RANGE			12:0
#define NVDLA_CDMA_D_DATAIN_SIZE_1_0_DATAIN_CHANNEL_SIZE				13


// Register NVDLA_CDMA_D_DATAIN_SIZE_EXT_0_0
#define NVDLA_CDMA_D_DATAIN_SIZE_EXT_0_0					32'h3024
#define NVDLA_CDMA_D_DATAIN_SIZE_EXT_0_0_DATAIN_WIDTH_EXT_RANGE			12:0
#define NVDLA_CDMA_D_DATAIN_SIZE_EXT_0_0_DATAIN_WIDTH_EXT_SIZE				13
#define NVDLA_CDMA_D_DATAIN_SIZE_EXT_0_0_DATAIN_HEIGHT_EXT_RANGE			28:16
#define NVDLA_CDMA_D_DATAIN_SIZE_EXT_0_0_DATAIN_HEIGHT_EXT_SIZE				13


// Register NVDLA_CDMA_D_PIXEL_OFFSET_0
#define NVDLA_CDMA_D_PIXEL_OFFSET_0					32'h3028
#define NVDLA_CDMA_D_PIXEL_OFFSET_0_PIXEL_X_OFFSET_RANGE			4:0
#define NVDLA_CDMA_D_PIXEL_OFFSET_0_PIXEL_X_OFFSET_SIZE				5
#define NVDLA_CDMA_D_PIXEL_OFFSET_0_PIXEL_Y_OFFSET_RANGE			18:16
#define NVDLA_CDMA_D_PIXEL_OFFSET_0_PIXEL_Y_OFFSET_SIZE				3


// Register NVDLA_CDMA_D_DAIN_RAM_TYPE_0
#define NVDLA_CDMA_D_DAIN_RAM_TYPE_0					32'h302c
#define NVDLA_CDMA_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_RANGE			0:0
#define NVDLA_CDMA_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_SIZE				1
#define NVDLA_CDMA_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_CVIF			1'h0
#define NVDLA_CDMA_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_MCIF			1'h1


// Register NVDLA_CDMA_D_DAIN_ADDR_HIGH_0_0
#define NVDLA_CDMA_D_DAIN_ADDR_HIGH_0_0					32'h3030
#define NVDLA_CDMA_D_DAIN_ADDR_HIGH_0_0_DATAIN_ADDR_HIGH_0_RANGE			31:0
#define NVDLA_CDMA_D_DAIN_ADDR_HIGH_0_0_DATAIN_ADDR_HIGH_0_SIZE				32


// Register NVDLA_CDMA_D_DAIN_ADDR_LOW_0_0
#define NVDLA_CDMA_D_DAIN_ADDR_LOW_0_0					32'h3034
#define NVDLA_CDMA_D_DAIN_ADDR_LOW_0_0_DATAIN_ADDR_LOW_0_RANGE			31:0
#define NVDLA_CDMA_D_DAIN_ADDR_LOW_0_0_DATAIN_ADDR_LOW_0_SIZE				32


// Register NVDLA_CDMA_D_DAIN_ADDR_HIGH_1_0
#define NVDLA_CDMA_D_DAIN_ADDR_HIGH_1_0					32'h3038
#define NVDLA_CDMA_D_DAIN_ADDR_HIGH_1_0_DATAIN_ADDR_HIGH_1_RANGE			31:0
#define NVDLA_CDMA_D_DAIN_ADDR_HIGH_1_0_DATAIN_ADDR_HIGH_1_SIZE				32


// Register NVDLA_CDMA_D_DAIN_ADDR_LOW_1_0
#define NVDLA_CDMA_D_DAIN_ADDR_LOW_1_0					32'h303c
#define NVDLA_CDMA_D_DAIN_ADDR_LOW_1_0_DATAIN_ADDR_LOW_1_RANGE			31:0
#define NVDLA_CDMA_D_DAIN_ADDR_LOW_1_0_DATAIN_ADDR_LOW_1_SIZE				32


// Register NVDLA_CDMA_D_LINE_STRIDE_0
#define NVDLA_CDMA_D_LINE_STRIDE_0					32'h3040
#define NVDLA_CDMA_D_LINE_STRIDE_0_LINE_STRIDE_RANGE			31:0
#define NVDLA_CDMA_D_LINE_STRIDE_0_LINE_STRIDE_SIZE				32


// Register NVDLA_CDMA_D_LINE_UV_STRIDE_0
#define NVDLA_CDMA_D_LINE_UV_STRIDE_0					32'h3044
#define NVDLA_CDMA_D_LINE_UV_STRIDE_0_UV_LINE_STRIDE_RANGE			31:0
#define NVDLA_CDMA_D_LINE_UV_STRIDE_0_UV_LINE_STRIDE_SIZE				32


// Register NVDLA_CDMA_D_SURF_STRIDE_0
#define NVDLA_CDMA_D_SURF_STRIDE_0					32'h3048
#define NVDLA_CDMA_D_SURF_STRIDE_0_SURF_STRIDE_RANGE			31:0
#define NVDLA_CDMA_D_SURF_STRIDE_0_SURF_STRIDE_SIZE				32


// Register NVDLA_CDMA_D_DAIN_MAP_0
#define NVDLA_CDMA_D_DAIN_MAP_0					32'h304c
#define NVDLA_CDMA_D_DAIN_MAP_0_LINE_PACKED_RANGE			0:0
#define NVDLA_CDMA_D_DAIN_MAP_0_LINE_PACKED_SIZE				1
#define NVDLA_CDMA_D_DAIN_MAP_0_LINE_PACKED_FALSE			1'h0
#define NVDLA_CDMA_D_DAIN_MAP_0_LINE_PACKED_TRUE			1'h1
#define NVDLA_CDMA_D_DAIN_MAP_0_SURF_PACKED_RANGE			16:16
#define NVDLA_CDMA_D_DAIN_MAP_0_SURF_PACKED_SIZE				1
#define NVDLA_CDMA_D_DAIN_MAP_0_SURF_PACKED_FALSE			1'h0
#define NVDLA_CDMA_D_DAIN_MAP_0_SURF_PACKED_TRUE			1'h1


// Register NVDLA_CDMA_D_RESERVED_X_CFG_0
#define NVDLA_CDMA_D_RESERVED_X_CFG_0					32'h3050
#define NVDLA_CDMA_D_RESERVED_X_CFG_0_RSV_PER_LINE_RANGE			9:0
#define NVDLA_CDMA_D_RESERVED_X_CFG_0_RSV_PER_LINE_SIZE				10
#define NVDLA_CDMA_D_RESERVED_X_CFG_0_RSV_PER_UV_LINE_RANGE			25:16
#define NVDLA_CDMA_D_RESERVED_X_CFG_0_RSV_PER_UV_LINE_SIZE				10


// Register NVDLA_CDMA_D_RESERVED_Y_CFG_0
#define NVDLA_CDMA_D_RESERVED_Y_CFG_0					32'h3054
#define NVDLA_CDMA_D_RESERVED_Y_CFG_0_RSV_HEIGHT_RANGE			2:0
#define NVDLA_CDMA_D_RESERVED_Y_CFG_0_RSV_HEIGHT_SIZE				3
#define NVDLA_CDMA_D_RESERVED_Y_CFG_0_RSV_Y_INDEX_RANGE			20:16
#define NVDLA_CDMA_D_RESERVED_Y_CFG_0_RSV_Y_INDEX_SIZE				5


// Register NVDLA_CDMA_D_BATCH_NUMBER_0
#define NVDLA_CDMA_D_BATCH_NUMBER_0					32'h3058
#define NVDLA_CDMA_D_BATCH_NUMBER_0_BATCHES_RANGE			4:0
#define NVDLA_CDMA_D_BATCH_NUMBER_0_BATCHES_SIZE				5


// Register NVDLA_CDMA_D_BATCH_STRIDE_0
#define NVDLA_CDMA_D_BATCH_STRIDE_0					32'h305c
#define NVDLA_CDMA_D_BATCH_STRIDE_0_BATCH_STRIDE_RANGE			31:0
#define NVDLA_CDMA_D_BATCH_STRIDE_0_BATCH_STRIDE_SIZE				32


// Register NVDLA_CDMA_D_ENTRY_PER_SLICE_0
#define NVDLA_CDMA_D_ENTRY_PER_SLICE_0					32'h3060
#define NVDLA_CDMA_D_ENTRY_PER_SLICE_0_ENTRIES_RANGE			13:0
#define NVDLA_CDMA_D_ENTRY_PER_SLICE_0_ENTRIES_SIZE				14


// Register NVDLA_CDMA_D_FETCH_GRAIN_0
#define NVDLA_CDMA_D_FETCH_GRAIN_0					32'h3064
#define NVDLA_CDMA_D_FETCH_GRAIN_0_GRAINS_RANGE			11:0
#define NVDLA_CDMA_D_FETCH_GRAIN_0_GRAINS_SIZE				12


// Register NVDLA_CDMA_D_WEIGHT_FORMAT_0
#define NVDLA_CDMA_D_WEIGHT_FORMAT_0					32'h3068
#define NVDLA_CDMA_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_RANGE			0:0
#define NVDLA_CDMA_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_SIZE				1
#define NVDLA_CDMA_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_UNCOMPRESSED			1'h0
#define NVDLA_CDMA_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_COMPRESSED			1'h1


// Register NVDLA_CDMA_D_WEIGHT_SIZE_0_0
#define NVDLA_CDMA_D_WEIGHT_SIZE_0_0					32'h306c
#define NVDLA_CDMA_D_WEIGHT_SIZE_0_0_BYTE_PER_KERNEL_RANGE			17:0
#define NVDLA_CDMA_D_WEIGHT_SIZE_0_0_BYTE_PER_KERNEL_SIZE				18


// Register NVDLA_CDMA_D_WEIGHT_SIZE_1_0
#define NVDLA_CDMA_D_WEIGHT_SIZE_1_0					32'h3070
#define NVDLA_CDMA_D_WEIGHT_SIZE_1_0_WEIGHT_KERNEL_RANGE			12:0
#define NVDLA_CDMA_D_WEIGHT_SIZE_1_0_WEIGHT_KERNEL_SIZE				13


// Register NVDLA_CDMA_D_WEIGHT_RAM_TYPE_0
#define NVDLA_CDMA_D_WEIGHT_RAM_TYPE_0					32'h3074
#define NVDLA_CDMA_D_WEIGHT_RAM_TYPE_0_WEIGHT_RAM_TYPE_RANGE			0:0
#define NVDLA_CDMA_D_WEIGHT_RAM_TYPE_0_WEIGHT_RAM_TYPE_SIZE				1
#define NVDLA_CDMA_D_WEIGHT_RAM_TYPE_0_WEIGHT_RAM_TYPE_CVIF			1'h0
#define NVDLA_CDMA_D_WEIGHT_RAM_TYPE_0_WEIGHT_RAM_TYPE_MCIF			1'h1


// Register NVDLA_CDMA_D_WEIGHT_ADDR_HIGH_0
#define NVDLA_CDMA_D_WEIGHT_ADDR_HIGH_0					32'h3078
#define NVDLA_CDMA_D_WEIGHT_ADDR_HIGH_0_WEIGHT_ADDR_HIGH_RANGE			31:0
#define NVDLA_CDMA_D_WEIGHT_ADDR_HIGH_0_WEIGHT_ADDR_HIGH_SIZE				32


// Register NVDLA_CDMA_D_WEIGHT_ADDR_LOW_0
#define NVDLA_CDMA_D_WEIGHT_ADDR_LOW_0					32'h307c
#define NVDLA_CDMA_D_WEIGHT_ADDR_LOW_0_WEIGHT_ADDR_LOW_RANGE			31:0
#define NVDLA_CDMA_D_WEIGHT_ADDR_LOW_0_WEIGHT_ADDR_LOW_SIZE				32


// Register NVDLA_CDMA_D_WEIGHT_BYTES_0
#define NVDLA_CDMA_D_WEIGHT_BYTES_0					32'h3080
#define NVDLA_CDMA_D_WEIGHT_BYTES_0_WEIGHT_BYTES_RANGE			31:0
#define NVDLA_CDMA_D_WEIGHT_BYTES_0_WEIGHT_BYTES_SIZE				32


// Register NVDLA_CDMA_D_WGS_ADDR_HIGH_0
#define NVDLA_CDMA_D_WGS_ADDR_HIGH_0					32'h3084
#define NVDLA_CDMA_D_WGS_ADDR_HIGH_0_WGS_ADDR_HIGH_RANGE			31:0
#define NVDLA_CDMA_D_WGS_ADDR_HIGH_0_WGS_ADDR_HIGH_SIZE				32


// Register NVDLA_CDMA_D_WGS_ADDR_LOW_0
#define NVDLA_CDMA_D_WGS_ADDR_LOW_0					32'h3088
#define NVDLA_CDMA_D_WGS_ADDR_LOW_0_WGS_ADDR_LOW_RANGE			31:0
#define NVDLA_CDMA_D_WGS_ADDR_LOW_0_WGS_ADDR_LOW_SIZE				32


// Register NVDLA_CDMA_D_WMB_ADDR_HIGH_0
#define NVDLA_CDMA_D_WMB_ADDR_HIGH_0					32'h308c
#define NVDLA_CDMA_D_WMB_ADDR_HIGH_0_WMB_ADDR_HIGH_RANGE			31:0
#define NVDLA_CDMA_D_WMB_ADDR_HIGH_0_WMB_ADDR_HIGH_SIZE				32


// Register NVDLA_CDMA_D_WMB_ADDR_LOW_0
#define NVDLA_CDMA_D_WMB_ADDR_LOW_0					32'h3090
#define NVDLA_CDMA_D_WMB_ADDR_LOW_0_WMB_ADDR_LOW_RANGE			31:0
#define NVDLA_CDMA_D_WMB_ADDR_LOW_0_WMB_ADDR_LOW_SIZE				32


// Register NVDLA_CDMA_D_WMB_BYTES_0
#define NVDLA_CDMA_D_WMB_BYTES_0					32'h3094
#define NVDLA_CDMA_D_WMB_BYTES_0_WMB_BYTES_RANGE			27:0
#define NVDLA_CDMA_D_WMB_BYTES_0_WMB_BYTES_SIZE				28


// Register NVDLA_CDMA_D_MEAN_FORMAT_0
#define NVDLA_CDMA_D_MEAN_FORMAT_0					32'h3098
#define NVDLA_CDMA_D_MEAN_FORMAT_0_MEAN_FORMAT_RANGE			0:0
#define NVDLA_CDMA_D_MEAN_FORMAT_0_MEAN_FORMAT_SIZE				1
#define NVDLA_CDMA_D_MEAN_FORMAT_0_MEAN_FORMAT_DISABLE			1'h0
#define NVDLA_CDMA_D_MEAN_FORMAT_0_MEAN_FORMAT_ENABLE			1'h1


// Register NVDLA_CDMA_D_MEAN_GLOBAL_0_0
#define NVDLA_CDMA_D_MEAN_GLOBAL_0_0					32'h309c
#define NVDLA_CDMA_D_MEAN_GLOBAL_0_0_MEAN_RY_RANGE			15:0
#define NVDLA_CDMA_D_MEAN_GLOBAL_0_0_MEAN_RY_SIZE				16
#define NVDLA_CDMA_D_MEAN_GLOBAL_0_0_MEAN_GU_RANGE			31:16
#define NVDLA_CDMA_D_MEAN_GLOBAL_0_0_MEAN_GU_SIZE				16


// Register NVDLA_CDMA_D_MEAN_GLOBAL_1_0
#define NVDLA_CDMA_D_MEAN_GLOBAL_1_0					32'h30a0
#define NVDLA_CDMA_D_MEAN_GLOBAL_1_0_MEAN_BV_RANGE			15:0
#define NVDLA_CDMA_D_MEAN_GLOBAL_1_0_MEAN_BV_SIZE				16
#define NVDLA_CDMA_D_MEAN_GLOBAL_1_0_MEAN_AX_RANGE			31:16
#define NVDLA_CDMA_D_MEAN_GLOBAL_1_0_MEAN_AX_SIZE				16


// Register NVDLA_CDMA_D_CVT_CFG_0
#define NVDLA_CDMA_D_CVT_CFG_0					32'h30a4
#define NVDLA_CDMA_D_CVT_CFG_0_CVT_EN_RANGE			0:0
#define NVDLA_CDMA_D_CVT_CFG_0_CVT_EN_SIZE				1
#define NVDLA_CDMA_D_CVT_CFG_0_CVT_EN_DISABLE			1'h0
#define NVDLA_CDMA_D_CVT_CFG_0_CVT_EN_ENABLE			1'h1
#define NVDLA_CDMA_D_CVT_CFG_0_CVT_TRUNCATE_RANGE			9:4
#define NVDLA_CDMA_D_CVT_CFG_0_CVT_TRUNCATE_SIZE				6


// Register NVDLA_CDMA_D_CVT_OFFSET_0
#define NVDLA_CDMA_D_CVT_OFFSET_0					32'h30a8
#define NVDLA_CDMA_D_CVT_OFFSET_0_CVT_OFFSET_RANGE			15:0
#define NVDLA_CDMA_D_CVT_OFFSET_0_CVT_OFFSET_SIZE				16


// Register NVDLA_CDMA_D_CVT_SCALE_0
#define NVDLA_CDMA_D_CVT_SCALE_0					32'h30ac
#define NVDLA_CDMA_D_CVT_SCALE_0_CVT_SCALE_RANGE			15:0
#define NVDLA_CDMA_D_CVT_SCALE_0_CVT_SCALE_SIZE				16


// Register NVDLA_CDMA_D_CONV_STRIDE_0
#define NVDLA_CDMA_D_CONV_STRIDE_0					32'h30b0
#define NVDLA_CDMA_D_CONV_STRIDE_0_CONV_X_STRIDE_RANGE			2:0
#define NVDLA_CDMA_D_CONV_STRIDE_0_CONV_X_STRIDE_SIZE				3
#define NVDLA_CDMA_D_CONV_STRIDE_0_CONV_Y_STRIDE_RANGE			18:16
#define NVDLA_CDMA_D_CONV_STRIDE_0_CONV_Y_STRIDE_SIZE				3


// Register NVDLA_CDMA_D_ZERO_PADDING_0
#define NVDLA_CDMA_D_ZERO_PADDING_0					32'h30b4
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_LEFT_RANGE			4:0
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_LEFT_SIZE				5
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_RIGHT_RANGE			13:8
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_RIGHT_SIZE				6
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_TOP_RANGE			20:16
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_TOP_SIZE				5
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_BOTTOM_RANGE			29:24
#define NVDLA_CDMA_D_ZERO_PADDING_0_PAD_BOTTOM_SIZE				6


// Register NVDLA_CDMA_D_ZERO_PADDING_VALUE_0
#define NVDLA_CDMA_D_ZERO_PADDING_VALUE_0					32'h30b8
#define NVDLA_CDMA_D_ZERO_PADDING_VALUE_0_PAD_VALUE_RANGE			15:0
#define NVDLA_CDMA_D_ZERO_PADDING_VALUE_0_PAD_VALUE_SIZE				16


// Register NVDLA_CDMA_D_BANK_0
#define NVDLA_CDMA_D_BANK_0					32'h30bc
#define NVDLA_CDMA_D_BANK_0_DATA_BANK_RANGE			4:0
#define NVDLA_CDMA_D_BANK_0_DATA_BANK_SIZE				5
#define NVDLA_CDMA_D_BANK_0_WEIGHT_BANK_RANGE			20:16
#define NVDLA_CDMA_D_BANK_0_WEIGHT_BANK_SIZE				5


// Register NVDLA_CDMA_D_NAN_FLUSH_TO_ZERO_0
#define NVDLA_CDMA_D_NAN_FLUSH_TO_ZERO_0					32'h30c0
#define NVDLA_CDMA_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_RANGE			0:0
#define NVDLA_CDMA_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_SIZE				1
#define NVDLA_CDMA_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_DISABLE			1'h0
#define NVDLA_CDMA_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_ENABLE			1'h1


// Register NVDLA_CDMA_D_NAN_INPUT_DATA_NUM_0
#define NVDLA_CDMA_D_NAN_INPUT_DATA_NUM_0					32'h30c4
#define NVDLA_CDMA_D_NAN_INPUT_DATA_NUM_0_NAN_DATA_NUM_RANGE			31:0
#define NVDLA_CDMA_D_NAN_INPUT_DATA_NUM_0_NAN_DATA_NUM_SIZE				32


// Register NVDLA_CDMA_D_NAN_INPUT_WEIGHT_NUM_0
#define NVDLA_CDMA_D_NAN_INPUT_WEIGHT_NUM_0					32'h30c8
#define NVDLA_CDMA_D_NAN_INPUT_WEIGHT_NUM_0_NAN_WEIGHT_NUM_RANGE			31:0
#define NVDLA_CDMA_D_NAN_INPUT_WEIGHT_NUM_0_NAN_WEIGHT_NUM_SIZE				32


// Register NVDLA_CDMA_D_INF_INPUT_DATA_NUM_0
#define NVDLA_CDMA_D_INF_INPUT_DATA_NUM_0					32'h30cc
#define NVDLA_CDMA_D_INF_INPUT_DATA_NUM_0_INF_DATA_NUM_RANGE			31:0
#define NVDLA_CDMA_D_INF_INPUT_DATA_NUM_0_INF_DATA_NUM_SIZE				32


// Register NVDLA_CDMA_D_INF_INPUT_WEIGHT_NUM_0
#define NVDLA_CDMA_D_INF_INPUT_WEIGHT_NUM_0					32'h30d0
#define NVDLA_CDMA_D_INF_INPUT_WEIGHT_NUM_0_INF_WEIGHT_NUM_RANGE			31:0
#define NVDLA_CDMA_D_INF_INPUT_WEIGHT_NUM_0_INF_WEIGHT_NUM_SIZE				32


// Register NVDLA_CDMA_D_PERF_ENABLE_0
#define NVDLA_CDMA_D_PERF_ENABLE_0					32'h30d4
#define NVDLA_CDMA_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_CDMA_D_PERF_ENABLE_0_DMA_EN_SIZE				1


// Register NVDLA_CDMA_D_PERF_DAT_READ_STALL_0
#define NVDLA_CDMA_D_PERF_DAT_READ_STALL_0					32'h30d8
#define NVDLA_CDMA_D_PERF_DAT_READ_STALL_0_DAT_RD_STALL_RANGE			31:0
#define NVDLA_CDMA_D_PERF_DAT_READ_STALL_0_DAT_RD_STALL_SIZE				32


// Register NVDLA_CDMA_D_PERF_WT_READ_STALL_0
#define NVDLA_CDMA_D_PERF_WT_READ_STALL_0					32'h30dc
#define NVDLA_CDMA_D_PERF_WT_READ_STALL_0_WT_RD_STALL_RANGE			31:0
#define NVDLA_CDMA_D_PERF_WT_READ_STALL_0_WT_RD_STALL_SIZE				32


// Register NVDLA_CDMA_D_PERF_DAT_READ_LATENCY_0
#define NVDLA_CDMA_D_PERF_DAT_READ_LATENCY_0					32'h30e0
#define NVDLA_CDMA_D_PERF_DAT_READ_LATENCY_0_DAT_RD_LATENCY_RANGE			31:0
#define NVDLA_CDMA_D_PERF_DAT_READ_LATENCY_0_DAT_RD_LATENCY_SIZE				32


// Register NVDLA_CDMA_D_PERF_WT_READ_LATENCY_0
#define NVDLA_CDMA_D_PERF_WT_READ_LATENCY_0					32'h30e4
#define NVDLA_CDMA_D_PERF_WT_READ_LATENCY_0_WT_RD_LATENCY_RANGE			31:0
#define NVDLA_CDMA_D_PERF_WT_READ_LATENCY_0_WT_RD_LATENCY_SIZE				32


// Register NVDLA_CDMA_D_CYA_0
#define NVDLA_CDMA_D_CYA_0					32'h30e8
#define NVDLA_CDMA_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CDMA_D_CYA_0_CYA_SIZE				32


// Register NVDLA_CSC_S_STATUS_0
#define NVDLA_CSC_S_STATUS_0					32'h4000
#define NVDLA_CSC_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CSC_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CSC_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CSC_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CSC_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CSC_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CSC_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CSC_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CSC_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CSC_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CSC_S_POINTER_0
#define NVDLA_CSC_S_POINTER_0					32'h4004
#define NVDLA_CSC_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CSC_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CSC_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CSC_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CSC_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CSC_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CSC_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CSC_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CSC_D_OP_ENABLE_0
#define NVDLA_CSC_D_OP_ENABLE_0					32'h4008
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CSC_D_MISC_CFG_0
#define NVDLA_CSC_D_MISC_CFG_0					32'h400c
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_RANGE			9:8
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_FP16			2'h2
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_RANGE			16:16
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_ENABLE			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_RANGE			20:20
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_ENABLE			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_RANGE			24:24
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_ENABLE			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_RANGE			28:28
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_ENABLE			1'h1


// Register NVDLA_CSC_D_DATAIN_FORMAT_0
#define NVDLA_CSC_D_DATAIN_FORMAT_0					32'h4010
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_RANGE			0:0
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_SIZE				1
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_FEATURE			1'h0
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_PIXEL			1'h1


// Register NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0					32'h4014
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_WIDTH_EXT_RANGE			12:0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_WIDTH_EXT_SIZE				13
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_HEIGHT_EXT_RANGE			28:16
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_HEIGHT_EXT_SIZE				13


// Register NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0					32'h4018
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0_DATAIN_CHANNEL_EXT_RANGE			12:0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0_DATAIN_CHANNEL_EXT_SIZE				13


// Register NVDLA_CSC_D_BATCH_NUMBER_0
#define NVDLA_CSC_D_BATCH_NUMBER_0					32'h401c
#define NVDLA_CSC_D_BATCH_NUMBER_0_BATCHES_RANGE			4:0
#define NVDLA_CSC_D_BATCH_NUMBER_0_BATCHES_SIZE				5


// Register NVDLA_CSC_D_POST_Y_EXTENSION_0
#define NVDLA_CSC_D_POST_Y_EXTENSION_0					32'h4020
#define NVDLA_CSC_D_POST_Y_EXTENSION_0_Y_EXTENSION_RANGE			1:0
#define NVDLA_CSC_D_POST_Y_EXTENSION_0_Y_EXTENSION_SIZE				2


// Register NVDLA_CSC_D_ENTRY_PER_SLICE_0
#define NVDLA_CSC_D_ENTRY_PER_SLICE_0					32'h4024
#define NVDLA_CSC_D_ENTRY_PER_SLICE_0_ENTRIES_RANGE			13:0
#define NVDLA_CSC_D_ENTRY_PER_SLICE_0_ENTRIES_SIZE				14


// Register NVDLA_CSC_D_WEIGHT_FORMAT_0
#define NVDLA_CSC_D_WEIGHT_FORMAT_0					32'h4028
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_RANGE			0:0
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_SIZE				1
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_UNCOMPRESSED			1'h0
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_COMPRESSED			1'h1


// Register NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0					32'h402c
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_WIDTH_EXT_RANGE			4:0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_WIDTH_EXT_SIZE				5
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_HEIGHT_EXT_RANGE			20:16
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_HEIGHT_EXT_SIZE				5


// Register NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0					32'h4030
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_CHANNEL_EXT_RANGE			12:0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_CHANNEL_EXT_SIZE				13
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_KERNEL_RANGE			28:16
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_KERNEL_SIZE				13


// Register NVDLA_CSC_D_WEIGHT_BYTES_0
#define NVDLA_CSC_D_WEIGHT_BYTES_0					32'h4034
#define NVDLA_CSC_D_WEIGHT_BYTES_0_WEIGHT_BYTES_RANGE			31:0
#define NVDLA_CSC_D_WEIGHT_BYTES_0_WEIGHT_BYTES_SIZE				32


// Register NVDLA_CSC_D_WMB_BYTES_0
#define NVDLA_CSC_D_WMB_BYTES_0					32'h4038
#define NVDLA_CSC_D_WMB_BYTES_0_WMB_BYTES_RANGE			27:0
#define NVDLA_CSC_D_WMB_BYTES_0_WMB_BYTES_SIZE				28


// Register NVDLA_CSC_D_DATAOUT_SIZE_0_0
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0					32'h403c
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_RANGE			12:0
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_SIZE				13
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_RANGE			28:16
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_SIZE				13


// Register NVDLA_CSC_D_DATAOUT_SIZE_1_0
#define NVDLA_CSC_D_DATAOUT_SIZE_1_0					32'h4040
#define NVDLA_CSC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_RANGE			12:0
#define NVDLA_CSC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_SIZE				13


// Register NVDLA_CSC_D_ATOMICS_0
#define NVDLA_CSC_D_ATOMICS_0					32'h4044
#define NVDLA_CSC_D_ATOMICS_0_ATOMICS_RANGE			20:0
#define NVDLA_CSC_D_ATOMICS_0_ATOMICS_SIZE				21


// Register NVDLA_CSC_D_RELEASE_0
#define NVDLA_CSC_D_RELEASE_0					32'h4048
#define NVDLA_CSC_D_RELEASE_0_RLS_SLICES_RANGE			11:0
#define NVDLA_CSC_D_RELEASE_0_RLS_SLICES_SIZE				12


// Register NVDLA_CSC_D_CONV_STRIDE_EXT_0
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0					32'h404c
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_X_STRIDE_EXT_RANGE			2:0
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_X_STRIDE_EXT_SIZE				3
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_Y_STRIDE_EXT_RANGE			18:16
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_Y_STRIDE_EXT_SIZE				3


// Register NVDLA_CSC_D_DILATION_EXT_0
#define NVDLA_CSC_D_DILATION_EXT_0					32'h4050
#define NVDLA_CSC_D_DILATION_EXT_0_X_DILATION_EXT_RANGE			4:0
#define NVDLA_CSC_D_DILATION_EXT_0_X_DILATION_EXT_SIZE				5
#define NVDLA_CSC_D_DILATION_EXT_0_Y_DILATION_EXT_RANGE			20:16
#define NVDLA_CSC_D_DILATION_EXT_0_Y_DILATION_EXT_SIZE				5


// Register NVDLA_CSC_D_ZERO_PADDING_0
#define NVDLA_CSC_D_ZERO_PADDING_0					32'h4054
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_LEFT_RANGE			4:0
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_LEFT_SIZE				5
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_TOP_RANGE			20:16
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_TOP_SIZE				5


// Register NVDLA_CSC_D_ZERO_PADDING_VALUE_0
#define NVDLA_CSC_D_ZERO_PADDING_VALUE_0					32'h4058
#define NVDLA_CSC_D_ZERO_PADDING_VALUE_0_PAD_VALUE_RANGE			15:0
#define NVDLA_CSC_D_ZERO_PADDING_VALUE_0_PAD_VALUE_SIZE				16


// Register NVDLA_CSC_D_BANK_0
#define NVDLA_CSC_D_BANK_0					32'h405c
#define NVDLA_CSC_D_BANK_0_DATA_BANK_RANGE			4:0
#define NVDLA_CSC_D_BANK_0_DATA_BANK_SIZE				5
#define NVDLA_CSC_D_BANK_0_WEIGHT_BANK_RANGE			20:16
#define NVDLA_CSC_D_BANK_0_WEIGHT_BANK_SIZE				5


// Register NVDLA_CSC_D_PRA_CFG_0
#define NVDLA_CSC_D_PRA_CFG_0					32'h4060
#define NVDLA_CSC_D_PRA_CFG_0_PRA_TRUNCATE_RANGE			1:0
#define NVDLA_CSC_D_PRA_CFG_0_PRA_TRUNCATE_SIZE				2


// Register NVDLA_CSC_D_CYA_0
#define NVDLA_CSC_D_CYA_0					32'h4064
#define NVDLA_CSC_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CSC_D_CYA_0_CYA_SIZE				32


// Register NVDLA_CMAC_A_S_STATUS_0
#define NVDLA_CMAC_A_S_STATUS_0					32'h5000
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CMAC_A_S_POINTER_0
#define NVDLA_CMAC_A_S_POINTER_0					32'h5004
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CMAC_A_D_OP_ENABLE_0
#define NVDLA_CMAC_A_D_OP_ENABLE_0					32'h5008
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CMAC_A_D_MISC_CFG_0
#define NVDLA_CMAC_A_D_MISC_CFG_0					32'h500c
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2


// Register NVDLA_CMAC_B_S_STATUS_0
#define NVDLA_CMAC_B_S_STATUS_0					32'h6000
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CMAC_B_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CMAC_B_S_POINTER_0
#define NVDLA_CMAC_B_S_POINTER_0					32'h6004
#define NVDLA_CMAC_B_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CMAC_B_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CMAC_B_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CMAC_B_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CMAC_B_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CMAC_B_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CMAC_B_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CMAC_B_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CMAC_B_D_OP_ENABLE_0
#define NVDLA_CMAC_B_D_OP_ENABLE_0					32'h6008
#define NVDLA_CMAC_B_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CMAC_B_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CMAC_B_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CMAC_B_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CMAC_B_D_MISC_CFG_0
#define NVDLA_CMAC_B_D_MISC_CFG_0					32'h600c
#define NVDLA_CMAC_B_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CMAC_B_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CMAC_B_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CMAC_B_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CMAC_B_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CMAC_B_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CMAC_B_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CMAC_B_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CMAC_B_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2


// Register NVDLA_CACC_S_STATUS_0
#define NVDLA_CACC_S_STATUS_0					32'h7000
#define NVDLA_CACC_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CACC_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CACC_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CACC_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CACC_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CACC_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CACC_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CACC_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CACC_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CACC_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CACC_S_POINTER_0
#define NVDLA_CACC_S_POINTER_0					32'h7004
#define NVDLA_CACC_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CACC_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CACC_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CACC_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CACC_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CACC_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CACC_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CACC_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CACC_D_OP_ENABLE_0
#define NVDLA_CACC_D_OP_ENABLE_0					32'h7008
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CACC_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CACC_D_MISC_CFG_0
#define NVDLA_CACC_D_MISC_CFG_0					32'h700c
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CACC_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CACC_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2


// Register NVDLA_CACC_D_DATAOUT_SIZE_0_0
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0					32'h7010
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_RANGE			12:0
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_SIZE				13
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_RANGE			28:16
#define NVDLA_CACC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_SIZE				13


// Register NVDLA_CACC_D_DATAOUT_SIZE_1_0
#define NVDLA_CACC_D_DATAOUT_SIZE_1_0					32'h7014
#define NVDLA_CACC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_RANGE			12:0
#define NVDLA_CACC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_SIZE				13


// Register NVDLA_CACC_D_DATAOUT_ADDR_0
#define NVDLA_CACC_D_DATAOUT_ADDR_0					32'h7018
#define NVDLA_CACC_D_DATAOUT_ADDR_0_DATAOUT_ADDR_RANGE			31:0
#define NVDLA_CACC_D_DATAOUT_ADDR_0_DATAOUT_ADDR_SIZE				32


// Register NVDLA_CACC_D_BATCH_NUMBER_0
#define NVDLA_CACC_D_BATCH_NUMBER_0					32'h701c
#define NVDLA_CACC_D_BATCH_NUMBER_0_BATCHES_RANGE			4:0
#define NVDLA_CACC_D_BATCH_NUMBER_0_BATCHES_SIZE				5


// Register NVDLA_CACC_D_LINE_STRIDE_0
#define NVDLA_CACC_D_LINE_STRIDE_0					32'h7020
#define NVDLA_CACC_D_LINE_STRIDE_0_LINE_STRIDE_RANGE			23:0
#define NVDLA_CACC_D_LINE_STRIDE_0_LINE_STRIDE_SIZE				24


// Register NVDLA_CACC_D_SURF_STRIDE_0
#define NVDLA_CACC_D_SURF_STRIDE_0					32'h7024
#define NVDLA_CACC_D_SURF_STRIDE_0_SURF_STRIDE_RANGE			23:0
#define NVDLA_CACC_D_SURF_STRIDE_0_SURF_STRIDE_SIZE				24


// Register NVDLA_CACC_D_DATAOUT_MAP_0
#define NVDLA_CACC_D_DATAOUT_MAP_0					32'h7028
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_RANGE			0:0
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_SIZE				1
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_FALSE			1'h0
#define NVDLA_CACC_D_DATAOUT_MAP_0_LINE_PACKED_TRUE			1'h1
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_RANGE			16:16
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_SIZE				1
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_FALSE			1'h0
#define NVDLA_CACC_D_DATAOUT_MAP_0_SURF_PACKED_TRUE			1'h1


// Register NVDLA_CACC_D_CLIP_CFG_0
#define NVDLA_CACC_D_CLIP_CFG_0					32'h702c
#define NVDLA_CACC_D_CLIP_CFG_0_CLIP_TRUNCATE_RANGE			4:0
#define NVDLA_CACC_D_CLIP_CFG_0_CLIP_TRUNCATE_SIZE				5


// Register NVDLA_CACC_D_OUT_SATURATION_0
#define NVDLA_CACC_D_OUT_SATURATION_0					32'h7030
#define NVDLA_CACC_D_OUT_SATURATION_0_SAT_COUNT_RANGE			31:0
#define NVDLA_CACC_D_OUT_SATURATION_0_SAT_COUNT_SIZE				32


// Register NVDLA_CACC_D_CYA_0
#define NVDLA_CACC_D_CYA_0					32'h7034
#define NVDLA_CACC_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CACC_D_CYA_0_CYA_SIZE				32


// Register NVDLA_SDP_RDMA_S_STATUS_0
#define NVDLA_SDP_RDMA_S_STATUS_0					32'h8000
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_SDP_RDMA_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_SDP_RDMA_S_POINTER_0
#define NVDLA_SDP_RDMA_S_POINTER_0					32'h8004
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_SDP_RDMA_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_SDP_RDMA_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_SDP_RDMA_D_OP_ENABLE_0
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0					32'h8008
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_SDP_RDMA_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0					32'h800c
#define NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0_WIDTH_RANGE			12:0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_WIDTH_0_WIDTH_SIZE				13


// Register NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0					32'h8010
#define NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0_HEIGHT_RANGE			12:0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_HEIGHT_0_HEIGHT_SIZE				13


// Register NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0					32'h8014
#define NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0_CHANNEL_RANGE			12:0
#define NVDLA_SDP_RDMA_D_DATA_CUBE_CHANNEL_0_CHANNEL_SIZE				13


// Register NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0					32'h8018
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0					32'h801c
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0					32'h8020
#define NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0					32'h8024
#define NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BRDMA_CFG_0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0					32'h8028
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_NO			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DISABLE_YES			1'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_RANGE			2:1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_SIZE				2
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_MUL			2'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_ALU			2'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_USE_BOTH			2'h2
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_RANGE			3:3
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_ONE_BYTE			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_SIZE_TWO_BYTE			1'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_RANGE			4:4
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_PER_KERNEL			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_DATA_MODE_PER_ELEMENT			1'h1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_RANGE			5:5
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_BRDMA_CFG_0_BRDMA_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0					32'h802c
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0_BS_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_LOW_0_BS_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0					32'h8030
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0_BS_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_BASE_ADDR_HIGH_0_BS_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0					32'h8034
#define NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0_BS_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_LINE_STRIDE_0_BS_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0					32'h8038
#define NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0_BS_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_SURFACE_STRIDE_0_BS_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0
#define NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0					32'h803c
#define NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0_BS_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BS_BATCH_STRIDE_0_BS_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_NRDMA_CFG_0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0					32'h8040
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_NO			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DISABLE_YES			1'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_RANGE			2:1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_SIZE				2
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_MUL			2'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_ALU			2'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_USE_BOTH			2'h2
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_RANGE			3:3
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_ONE_BYTE			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_SIZE_TWO_BYTE			1'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_RANGE			4:4
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_PER_KERNEL			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_DATA_MODE_PER_ELEMENT			1'h1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_RANGE			5:5
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_NRDMA_CFG_0_NRDMA_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0					32'h8044
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0_BN_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_LOW_0_BN_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0					32'h8048
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0_BN_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_BASE_ADDR_HIGH_0_BN_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0					32'h804c
#define NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0_BN_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_LINE_STRIDE_0_BN_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0					32'h8050
#define NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0_BN_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_SURFACE_STRIDE_0_BN_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0
#define NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0					32'h8054
#define NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0_BN_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_BN_BATCH_STRIDE_0_BN_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_ERDMA_CFG_0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0					32'h8058
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_NO			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DISABLE_YES			1'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_RANGE			2:1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_SIZE				2
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_MUL			2'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_ALU			2'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_USE_BOTH			2'h2
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_RANGE			3:3
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_ONE_BYTE			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_SIZE_TWO_BYTE			1'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_RANGE			4:4
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_PER_KERNEL			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_DATA_MODE_PER_ELEMENT			1'h1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_RANGE			5:5
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_ERDMA_CFG_0_ERDMA_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0					32'h805c
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0_EW_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_LOW_0_EW_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0					32'h8060
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0_EW_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_BASE_ADDR_HIGH_0_EW_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0
#define NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0					32'h8064
#define NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0_EW_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_LINE_STRIDE_0_EW_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0
#define NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0					32'h8068
#define NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0_EW_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_SURFACE_STRIDE_0_EW_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0
#define NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0					32'h806c
#define NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0_EW_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_RDMA_D_EW_BATCH_STRIDE_0_EW_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0					32'h8070
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_SIZE				1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_OFF			1'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_FLYING_MODE_ON			1'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_RANGE			1:1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_SIZE				1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_OFF			1'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_WINOGRAD_ON			1'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_RANGE			3:2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_IN_PRECISION_FP16			2'h2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_RANGE			5:4
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_RANGE			7:6
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_SIZE				2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_INT8			2'h0
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_INT16			2'h1
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_OUT_PRECISION_FP16			2'h2
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_RANGE			12:8
#define NVDLA_SDP_RDMA_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_SIZE				5


// Register NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0					32'h8074
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_RANGE			0:0
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_SIZE				1
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0
#define NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0					32'h8078
#define NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_RDMA_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0
#define NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0					32'h807c
#define NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_RDMA_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_ENABLE_0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0					32'h8080
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_RANGE			0:0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_SIZE				1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_NO			1'h0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_DMA_EN_YES			1'h1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_RANGE			1:1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_SIZE				1
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_NO			1'h0
#define NVDLA_SDP_RDMA_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_YES			1'h1


// Register NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0					32'h8084
#define NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0_MRDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_MRDMA_READ_STALL_0_MRDMA_STALL_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0					32'h8088
#define NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0_BRDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_BRDMA_READ_STALL_0_BRDMA_STALL_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0					32'h808c
#define NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0_NRDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_NRDMA_READ_STALL_0_NRDMA_STALL_SIZE				32


// Register NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0
#define NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0					32'h8090
#define NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0_ERDMA_STALL_RANGE			31:0
#define NVDLA_SDP_RDMA_D_PERF_ERDMA_READ_STALL_0_ERDMA_STALL_SIZE				32


// Register NVDLA_SDP_S_STATUS_0
#define NVDLA_SDP_S_STATUS_0					32'h9000
#define NVDLA_SDP_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_SDP_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_SDP_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_SDP_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_SDP_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_SDP_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_SDP_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_SDP_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_SDP_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_SDP_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_SDP_S_POINTER_0
#define NVDLA_SDP_S_POINTER_0					32'h9004
#define NVDLA_SDP_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_SDP_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_SDP_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_SDP_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_SDP_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_SDP_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_SDP_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_SDP_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_SDP_S_LUT_ACCESS_CFG_0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0					32'h9008
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ADDR_RANGE			9:0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ADDR_SIZE				10
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_RANGE			16:16
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_SIZE				1
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_LE			1'h0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_LO			1'h1
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_RANGE			17:17
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_SIZE				1
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_READ			1'h0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_WRITE			1'h1


// Register NVDLA_SDP_S_LUT_ACCESS_DATA_0
#define NVDLA_SDP_S_LUT_ACCESS_DATA_0					32'h900c
#define NVDLA_SDP_S_LUT_ACCESS_DATA_0_LUT_DATA_RANGE			15:0
#define NVDLA_SDP_S_LUT_ACCESS_DATA_0_LUT_DATA_SIZE				16


// Register NVDLA_SDP_S_LUT_CFG_0
#define NVDLA_SDP_S_LUT_CFG_0					32'h9010
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_RANGE			0:0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_EXPONENT			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_LINEAR			1'h1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_RANGE			4:4
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_LE			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_LO			1'h1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_RANGE			5:5
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_LE			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_LO			1'h1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_RANGE			6:6
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_LE			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_LO			1'h1


// Register NVDLA_SDP_S_LUT_INFO_0
#define NVDLA_SDP_S_LUT_INFO_0					32'h9014
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_OFFSET_RANGE			7:0
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_OFFSET_SIZE				8
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_SELECT_RANGE			15:8
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_SELECT_SIZE				8
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LO_INDEX_SELECT_RANGE			23:16
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LO_INDEX_SELECT_SIZE				8


// Register NVDLA_SDP_S_LUT_LE_START_0
#define NVDLA_SDP_S_LUT_LE_START_0					32'h9018
#define NVDLA_SDP_S_LUT_LE_START_0_LUT_LE_START_RANGE			31:0
#define NVDLA_SDP_S_LUT_LE_START_0_LUT_LE_START_SIZE				32


// Register NVDLA_SDP_S_LUT_LE_END_0
#define NVDLA_SDP_S_LUT_LE_END_0					32'h901c
#define NVDLA_SDP_S_LUT_LE_END_0_LUT_LE_END_RANGE			31:0
#define NVDLA_SDP_S_LUT_LE_END_0_LUT_LE_END_SIZE				32


// Register NVDLA_SDP_S_LUT_LO_START_0
#define NVDLA_SDP_S_LUT_LO_START_0					32'h9020
#define NVDLA_SDP_S_LUT_LO_START_0_LUT_LO_START_RANGE			31:0
#define NVDLA_SDP_S_LUT_LO_START_0_LUT_LO_START_SIZE				32


// Register NVDLA_SDP_S_LUT_LO_END_0
#define NVDLA_SDP_S_LUT_LO_END_0					32'h9024
#define NVDLA_SDP_S_LUT_LO_END_0_LUT_LO_END_RANGE			31:0
#define NVDLA_SDP_S_LUT_LO_END_0_LUT_LO_END_SIZE				32


// Register NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0					32'h9028
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_UFLOW_SCALE_RANGE			15:0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_UFLOW_SCALE_SIZE				16
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_OFLOW_SCALE_RANGE			31:16
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_OFLOW_SCALE_SIZE				16


// Register NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0					32'h902c
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_UFLOW_SHIFT_RANGE			4:0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_UFLOW_SHIFT_SIZE				5
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_OFLOW_SHIFT_RANGE			9:5
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_OFLOW_SHIFT_SIZE				5


// Register NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0					32'h9030
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_UFLOW_SCALE_RANGE			15:0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_UFLOW_SCALE_SIZE				16
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_OFLOW_SCALE_RANGE			31:16
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_OFLOW_SCALE_SIZE				16


// Register NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0					32'h9034
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_UFLOW_SHIFT_RANGE			4:0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_UFLOW_SHIFT_SIZE				5
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_OFLOW_SHIFT_RANGE			9:5
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_OFLOW_SHIFT_SIZE				5


// Register NVDLA_SDP_D_OP_ENABLE_0
#define NVDLA_SDP_D_OP_ENABLE_0					32'h9038
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_SDP_D_DATA_CUBE_WIDTH_0
#define NVDLA_SDP_D_DATA_CUBE_WIDTH_0					32'h903c
#define NVDLA_SDP_D_DATA_CUBE_WIDTH_0_WIDTH_RANGE			12:0
#define NVDLA_SDP_D_DATA_CUBE_WIDTH_0_WIDTH_SIZE				13


// Register NVDLA_SDP_D_DATA_CUBE_HEIGHT_0
#define NVDLA_SDP_D_DATA_CUBE_HEIGHT_0					32'h9040
#define NVDLA_SDP_D_DATA_CUBE_HEIGHT_0_HEIGHT_RANGE			12:0
#define NVDLA_SDP_D_DATA_CUBE_HEIGHT_0_HEIGHT_SIZE				13


// Register NVDLA_SDP_D_DATA_CUBE_CHANNEL_0
#define NVDLA_SDP_D_DATA_CUBE_CHANNEL_0					32'h9044
#define NVDLA_SDP_D_DATA_CUBE_CHANNEL_0_CHANNEL_RANGE			12:0
#define NVDLA_SDP_D_DATA_CUBE_CHANNEL_0_CHANNEL_SIZE				13


// Register NVDLA_SDP_D_DST_BASE_ADDR_LOW_0
#define NVDLA_SDP_D_DST_BASE_ADDR_LOW_0					32'h9048
#define NVDLA_SDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0
#define NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0					32'h904c
#define NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_D_DST_LINE_STRIDE_0
#define NVDLA_SDP_D_DST_LINE_STRIDE_0					32'h9050
#define NVDLA_SDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_D_DST_SURFACE_STRIDE_0
#define NVDLA_SDP_D_DST_SURFACE_STRIDE_0					32'h9054
#define NVDLA_SDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_D_DP_BS_CFG_0
#define NVDLA_SDP_D_DP_BS_CFG_0					32'h9058
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_RANGE			0:0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_RANGE			3:2
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_SIZE				2
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_MAX			2'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_MIN			2'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_SUM			2'h2
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_RANGE			4:4
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_RANGE			5:5
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_RANGE			6:6
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_BS_ALU_CFG_0
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0					32'h905c
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SHIFT_VALUE_RANGE			13:8
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SHIFT_VALUE_SIZE				6


// Register NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0					32'h9060
#define NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0_BS_ALU_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0_BS_ALU_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_BS_MUL_CFG_0
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0					32'h9064
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SHIFT_VALUE_RANGE			15:8
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SHIFT_VALUE_SIZE				8


// Register NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0					32'h9068
#define NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0_BS_MUL_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0_BS_MUL_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_BN_CFG_0
#define NVDLA_SDP_D_DP_BN_CFG_0					32'h906c
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_RANGE			0:0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_RANGE			3:2
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_SIZE				2
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_MAX			2'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_MIN			2'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_SUM			2'h2
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_RANGE			4:4
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_RANGE			5:5
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_RANGE			6:6
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_BN_ALU_CFG_0
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0					32'h9070
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SHIFT_VALUE_RANGE			13:8
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SHIFT_VALUE_SIZE				6


// Register NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0					32'h9074
#define NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0_BN_ALU_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0_BN_ALU_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_BN_MUL_CFG_0
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0					32'h9078
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SHIFT_VALUE_RANGE			15:8
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SHIFT_VALUE_SIZE				8


// Register NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0					32'h907c
#define NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0_BN_MUL_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0_BN_MUL_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_EW_CFG_0
#define NVDLA_SDP_D_DP_EW_CFG_0					32'h9080
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_RANGE			0:0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_RANGE			3:2
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_SIZE				2
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_MAX			2'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_MIN			2'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_SUM			2'h2
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_EQL			2'h3
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_RANGE			4:4
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_RANGE			5:5
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_RANGE			6:6
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_EW_ALU_CFG_0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0					32'h9084
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_SIZE				1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0					32'h9088
#define NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0_EW_ALU_OPERAND_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0_EW_ALU_OPERAND_SIZE				32


// Register NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0					32'h908c
#define NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0_EW_ALU_CVT_OFFSET_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0_EW_ALU_CVT_OFFSET_SIZE				32


// Register NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0					32'h9090
#define NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0_EW_ALU_CVT_SCALE_RANGE			15:0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0_EW_ALU_CVT_SCALE_SIZE				16


// Register NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0					32'h9094
#define NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0_EW_ALU_CVT_TRUNCATE_RANGE			5:0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0_EW_ALU_CVT_TRUNCATE_SIZE				6


// Register NVDLA_SDP_D_DP_EW_MUL_CFG_0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0					32'h9098
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_SIZE				1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0					32'h909c
#define NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0_EW_MUL_OPERAND_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0_EW_MUL_OPERAND_SIZE				32


// Register NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0					32'h90a0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0_EW_MUL_CVT_OFFSET_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0_EW_MUL_CVT_OFFSET_SIZE				32


// Register NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0					32'h90a4
#define NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0_EW_MUL_CVT_SCALE_RANGE			15:0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0_EW_MUL_CVT_SCALE_SIZE				16


// Register NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0					32'h90a8
#define NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0_EW_MUL_CVT_TRUNCATE_RANGE			5:0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0_EW_MUL_CVT_TRUNCATE_SIZE				6


// Register NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0
#define NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0					32'h90ac
#define NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0_EW_TRUNCATE_RANGE			9:0
#define NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0_EW_TRUNCATE_SIZE				10


// Register NVDLA_SDP_D_FEATURE_MODE_CFG_0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0					32'h90b0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_RANGE			0:0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_OFF			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_ON			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_RANGE			1:1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_MEM			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_PDP			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_RANGE			2:2
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_OFF			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_ON			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_RANGE			3:3
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_DISABLE			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_ENABLE			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_RANGE			12:8
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_SIZE				5


// Register NVDLA_SDP_D_DST_DMA_CFG_0
#define NVDLA_SDP_D_DST_DMA_CFG_0					32'h90b4
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_RANGE			0:0
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_SIZE				1
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_D_DST_BATCH_STRIDE_0
#define NVDLA_SDP_D_DST_BATCH_STRIDE_0					32'h90b8
#define NVDLA_SDP_D_DST_BATCH_STRIDE_0_DST_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_D_DST_BATCH_STRIDE_0_DST_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_D_DATA_FORMAT_0
#define NVDLA_SDP_D_DATA_FORMAT_0					32'h90bc
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_RANGE			1:0
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_SIZE				2
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_RANGE			3:2
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_SIZE				2
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_INT8			2'h0
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_INT16			2'h1
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_FP16			2'h2


// Register NVDLA_SDP_D_CVT_OFFSET_0
#define NVDLA_SDP_D_CVT_OFFSET_0					32'h90c0
#define NVDLA_SDP_D_CVT_OFFSET_0_CVT_OFFSET_RANGE			31:0
#define NVDLA_SDP_D_CVT_OFFSET_0_CVT_OFFSET_SIZE				32


// Register NVDLA_SDP_D_CVT_SCALE_0
#define NVDLA_SDP_D_CVT_SCALE_0					32'h90c4
#define NVDLA_SDP_D_CVT_SCALE_0_CVT_SCALE_RANGE			15:0
#define NVDLA_SDP_D_CVT_SCALE_0_CVT_SCALE_SIZE				16


// Register NVDLA_SDP_D_CVT_SHIFT_0
#define NVDLA_SDP_D_CVT_SHIFT_0					32'h90c8
#define NVDLA_SDP_D_CVT_SHIFT_0_CVT_SHIFT_RANGE			5:0
#define NVDLA_SDP_D_CVT_SHIFT_0_CVT_SHIFT_SIZE				6


// Register NVDLA_SDP_D_STATUS_0
#define NVDLA_SDP_D_STATUS_0					32'h90cc
#define NVDLA_SDP_D_STATUS_0_STATUS_UNEQUAL_RANGE			0:0
#define NVDLA_SDP_D_STATUS_0_STATUS_UNEQUAL_SIZE				1


// Register NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0
#define NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0					32'h90d0
#define NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0
#define NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0					32'h90d4
#define NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0
#define NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0					32'h90d8
#define NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0_STATUS_NAN_OUTPUT_NUM_RANGE			31:0
#define NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0_STATUS_NAN_OUTPUT_NUM_SIZE				32


// Register NVDLA_SDP_D_PERF_ENABLE_0
#define NVDLA_SDP_D_PERF_ENABLE_0					32'h90dc
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_RANGE			0:0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_YES			1'h1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_RANGE			1:1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_YES			1'h1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_RANGE			2:2
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_YES			1'h1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_RANGE			3:3
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_YES			1'h1


// Register NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0
#define NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0					32'h90e0
#define NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0_WDMA_STALL_RANGE			31:0
#define NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0_WDMA_STALL_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_UFLOW_0
#define NVDLA_SDP_D_PERF_LUT_UFLOW_0					32'h90e4
#define NVDLA_SDP_D_PERF_LUT_UFLOW_0_LUT_UFLOW_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_UFLOW_0_LUT_UFLOW_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_OFLOW_0
#define NVDLA_SDP_D_PERF_LUT_OFLOW_0					32'h90e8
#define NVDLA_SDP_D_PERF_LUT_OFLOW_0_LUT_OFLOW_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_OFLOW_0_LUT_OFLOW_SIZE				32


// Register NVDLA_SDP_D_PERF_OUT_SATURATION_0
#define NVDLA_SDP_D_PERF_OUT_SATURATION_0					32'h90ec
#define NVDLA_SDP_D_PERF_OUT_SATURATION_0_OUT_SATURATION_RANGE			31:0
#define NVDLA_SDP_D_PERF_OUT_SATURATION_0_OUT_SATURATION_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_HYBRID_0
#define NVDLA_SDP_D_PERF_LUT_HYBRID_0					32'h90f0
#define NVDLA_SDP_D_PERF_LUT_HYBRID_0_LUT_HYBRID_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_HYBRID_0_LUT_HYBRID_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_LE_HIT_0
#define NVDLA_SDP_D_PERF_LUT_LE_HIT_0					32'h90f4
#define NVDLA_SDP_D_PERF_LUT_LE_HIT_0_LUT_LE_HIT_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_LE_HIT_0_LUT_LE_HIT_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_LO_HIT_0
#define NVDLA_SDP_D_PERF_LUT_LO_HIT_0					32'h90f8
#define NVDLA_SDP_D_PERF_LUT_LO_HIT_0_LUT_LO_HIT_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_LO_HIT_0_LUT_LO_HIT_SIZE				32


// Register NVDLA_PDP_RDMA_S_STATUS_0
#define NVDLA_PDP_RDMA_S_STATUS_0					32'ha000
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_PDP_RDMA_S_POINTER_0
#define NVDLA_PDP_RDMA_S_POINTER_0					32'ha004
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_PDP_RDMA_D_OP_ENABLE_0
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0					32'ha008
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0					32'ha00c
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_RANGE			12:0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_SIZE				13


// Register NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0					32'ha010
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_RANGE			12:0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_SIZE				13


// Register NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0					32'ha014
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_RANGE			12:0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_SIZE				13


// Register NVDLA_PDP_RDMA_D_FLYING_MODE_0
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0					32'ha018
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_RANGE			0:0
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_SIZE				1
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_ON_FLYING			1'h0
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_OFF_FLYING			1'h1


// Register NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0					32'ha01c
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0					32'ha020
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0
#define NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0					32'ha024
#define NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0
#define NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0					32'ha028
#define NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0					32'ha02c
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_RANGE			0:0
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_SIZE				1
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_CV			1'h0
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_MC			1'h1


// Register NVDLA_PDP_RDMA_D_DATA_FORMAT_0
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0					32'ha030
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_RANGE			1:0
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_SIZE				2
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_INT8			2'h0
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_INT16			2'h1
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_FP16			2'h2


// Register NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0
#define NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0					32'ha034
#define NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0_SPLIT_NUM_RANGE			7:0
#define NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0_SPLIT_NUM_SIZE				8


// Register NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0					32'ha038
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_RANGE			3:0
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_SIZE				4
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_1			4'h0
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_2			4'h1
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_3			4'h2
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_4			4'h3
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_5			4'h4
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_6			4'h5
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_7			4'h6
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_8			4'h7
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_RANGE			7:4
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_SIZE				4


// Register NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0
#define NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0					32'ha03c
#define NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0_PAD_WIDTH_RANGE			3:0
#define NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0_PAD_WIDTH_SIZE				4


// Register NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0					32'ha040
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_RANGE			9:0
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_SIZE				10
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_RANGE			19:10
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_SIZE				10
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_RANGE			29:20
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_SIZE				10


// Register NVDLA_PDP_RDMA_D_PERF_ENABLE_0
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0					32'ha044
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_SIZE				1
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_DISABLE			1'h0
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_ENABLE			1'h1


// Register NVDLA_PDP_RDMA_D_PERF_READ_STALL_0
#define NVDLA_PDP_RDMA_D_PERF_READ_STALL_0					32'ha048
#define NVDLA_PDP_RDMA_D_PERF_READ_STALL_0_PERF_READ_STALL_RANGE			31:0
#define NVDLA_PDP_RDMA_D_PERF_READ_STALL_0_PERF_READ_STALL_SIZE				32


// Register NVDLA_PDP_RDMA_D_CYA_0
#define NVDLA_PDP_RDMA_D_CYA_0					32'ha04c
#define NVDLA_PDP_RDMA_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_PDP_RDMA_D_CYA_0_CYA_SIZE				32


// Register NVDLA_PDP_S_STATUS_0
#define NVDLA_PDP_S_STATUS_0					32'hb000
#define NVDLA_PDP_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_PDP_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_PDP_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_PDP_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_PDP_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_PDP_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_PDP_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_PDP_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_PDP_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_PDP_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_PDP_S_POINTER_0
#define NVDLA_PDP_S_POINTER_0					32'hb004
#define NVDLA_PDP_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_PDP_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_PDP_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_PDP_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_PDP_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_PDP_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_PDP_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_PDP_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_PDP_D_OP_ENABLE_0
#define NVDLA_PDP_D_OP_ENABLE_0					32'hb008
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_PDP_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0
#define NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0					32'hb00c
#define NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0
#define NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0					32'hb010
#define NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0
#define NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0					32'hb014
#define NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0
#define NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0					32'hb018
#define NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0_CUBE_OUT_WIDTH_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_OUT_WIDTH_0_CUBE_OUT_WIDTH_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0
#define NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0					32'hb01c
#define NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0_CUBE_OUT_HEIGHT_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_OUT_HEIGHT_0_CUBE_OUT_HEIGHT_SIZE				13


// Register NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0
#define NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0					32'hb020
#define NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0_CUBE_OUT_CHANNEL_RANGE			12:0
#define NVDLA_PDP_D_DATA_CUBE_OUT_CHANNEL_0_CUBE_OUT_CHANNEL_SIZE				13


// Register NVDLA_PDP_D_OPERATION_MODE_CFG_0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0					32'hb024
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_RANGE			1:0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_SIZE				2
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_POOLING_METHOD_AVERAGE			2'h0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_POOLING_METHOD_MAX			2'h1
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_POOLING_METHOD_POOLING_METHOD_MIN			2'h2
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_RANGE			4:4
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_SIZE				1
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_ON_FLYING			1'h0
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_FLYING_MODE_OFF_FLYING			1'h1
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_SPLIT_NUM_RANGE			15:8
#define NVDLA_PDP_D_OPERATION_MODE_CFG_0_SPLIT_NUM_SIZE				8


// Register NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0					32'hb028
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_RANGE			0:0
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_SIZE				1
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_DISABLE			1'h0
#define NVDLA_PDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_ENABLE			1'h1


// Register NVDLA_PDP_D_PARTIAL_WIDTH_IN_0
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0					32'hb02c
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_RANGE			9:0
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_RANGE			19:10
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_RANGE			29:20
#define NVDLA_PDP_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_SIZE				10


// Register NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0					32'hb030
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_FIRST_RANGE			9:0
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_FIRST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_LAST_RANGE			19:10
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_LAST_SIZE				10
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_MID_RANGE			29:20
#define NVDLA_PDP_D_PARTIAL_WIDTH_OUT_0_PARTIAL_WIDTH_OUT_MID_SIZE				10


// Register NVDLA_PDP_D_POOLING_KERNEL_CFG_0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0					32'hb034
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_RANGE			3:0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_SIZE				4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_1			4'h0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_2			4'h1
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_3			4'h2
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_4			4'h3
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_5			4'h4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_6			4'h5
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_7			4'h6
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_8			4'h7
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_RANGE			11:8
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_SIZE				4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_1			4'h0
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_2			4'h1
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_3			4'h2
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_4			4'h3
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_5			4'h4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_6			4'h5
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_7			4'h6
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_HEIGHT_KERNEL_HEIGHT_8			4'h7
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_RANGE			19:16
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_SIZE				4
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_HEIGHT_RANGE			23:20
#define NVDLA_PDP_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_HEIGHT_SIZE				4


// Register NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0
#define NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0					32'hb038
#define NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0_RECIP_KERNEL_WIDTH_RANGE			16:0
#define NVDLA_PDP_D_RECIP_KERNEL_WIDTH_0_RECIP_KERNEL_WIDTH_SIZE				17


// Register NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0
#define NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0					32'hb03c
#define NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0_RECIP_KERNEL_HEIGHT_RANGE			16:0
#define NVDLA_PDP_D_RECIP_KERNEL_HEIGHT_0_RECIP_KERNEL_HEIGHT_SIZE				17


// Register NVDLA_PDP_D_POOLING_PADDING_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0					32'hb040
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_LEFT_RANGE			2:0
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_LEFT_SIZE				3
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_TOP_RANGE			6:4
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_TOP_SIZE				3
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_RIGHT_RANGE			10:8
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_RIGHT_SIZE				3
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_BOTTOM_RANGE			14:12
#define NVDLA_PDP_D_POOLING_PADDING_CFG_0_PAD_BOTTOM_SIZE				3


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0					32'hb044
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0_PAD_VALUE_1X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_1_CFG_0_PAD_VALUE_1X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0					32'hb048
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0_PAD_VALUE_2X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_2_CFG_0_PAD_VALUE_2X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0					32'hb04c
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0_PAD_VALUE_3X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_3_CFG_0_PAD_VALUE_3X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0					32'hb050
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0_PAD_VALUE_4X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_4_CFG_0_PAD_VALUE_4X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0					32'hb054
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0_PAD_VALUE_5X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_5_CFG_0_PAD_VALUE_5X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0					32'hb058
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0_PAD_VALUE_6X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_6_CFG_0_PAD_VALUE_6X_SIZE				19


// Register NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0					32'hb05c
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0_PAD_VALUE_7X_RANGE			18:0
#define NVDLA_PDP_D_POOLING_PADDING_VALUE_7_CFG_0_PAD_VALUE_7X_SIZE				19


// Register NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0					32'hb060
#define NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_PDP_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0					32'hb064
#define NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_PDP_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_PDP_D_SRC_LINE_STRIDE_0
#define NVDLA_PDP_D_SRC_LINE_STRIDE_0					32'hb068
#define NVDLA_PDP_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_SRC_SURFACE_STRIDE_0
#define NVDLA_PDP_D_SRC_SURFACE_STRIDE_0					32'hb06c
#define NVDLA_PDP_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_DST_BASE_ADDR_LOW_0
#define NVDLA_PDP_D_DST_BASE_ADDR_LOW_0					32'hb070
#define NVDLA_PDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_PDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0
#define NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0					32'hb074
#define NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_PDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_PDP_D_DST_LINE_STRIDE_0
#define NVDLA_PDP_D_DST_LINE_STRIDE_0					32'hb078
#define NVDLA_PDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_DST_SURFACE_STRIDE_0
#define NVDLA_PDP_D_DST_SURFACE_STRIDE_0					32'hb07c
#define NVDLA_PDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_PDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_SIZE				32


// Register NVDLA_PDP_D_DST_RAM_CFG_0
#define NVDLA_PDP_D_DST_RAM_CFG_0					32'hb080
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_RANGE			0:0
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_SIZE				1
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_CV			1'h0
#define NVDLA_PDP_D_DST_RAM_CFG_0_DST_RAM_TYPE_MC			1'h1


// Register NVDLA_PDP_D_DATA_FORMAT_0
#define NVDLA_PDP_D_DATA_FORMAT_0					32'hb084
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_RANGE			1:0
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_SIZE				2
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_INT8			2'h0
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_INT16			2'h1
#define NVDLA_PDP_D_DATA_FORMAT_0_INPUT_DATA_FP16			2'h2


// Register NVDLA_PDP_D_INF_INPUT_NUM_0
#define NVDLA_PDP_D_INF_INPUT_NUM_0					32'hb088
#define NVDLA_PDP_D_INF_INPUT_NUM_0_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_PDP_D_INF_INPUT_NUM_0_INF_INPUT_NUM_SIZE				32


// Register NVDLA_PDP_D_NAN_INPUT_NUM_0
#define NVDLA_PDP_D_NAN_INPUT_NUM_0					32'hb08c
#define NVDLA_PDP_D_NAN_INPUT_NUM_0_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_PDP_D_NAN_INPUT_NUM_0_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_PDP_D_NAN_OUTPUT_NUM_0
#define NVDLA_PDP_D_NAN_OUTPUT_NUM_0					32'hb090
#define NVDLA_PDP_D_NAN_OUTPUT_NUM_0_NAN_OUTPUT_NUM_RANGE			31:0
#define NVDLA_PDP_D_NAN_OUTPUT_NUM_0_NAN_OUTPUT_NUM_SIZE				32


// Register NVDLA_PDP_D_PERF_ENABLE_0
#define NVDLA_PDP_D_PERF_ENABLE_0					32'hb094
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_SIZE				1
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_DISABLE			1'h0
#define NVDLA_PDP_D_PERF_ENABLE_0_DMA_EN_ENABLE			1'h1


// Register NVDLA_PDP_D_PERF_WRITE_STALL_0
#define NVDLA_PDP_D_PERF_WRITE_STALL_0					32'hb098
#define NVDLA_PDP_D_PERF_WRITE_STALL_0_PERF_WRITE_STALL_RANGE			31:0
#define NVDLA_PDP_D_PERF_WRITE_STALL_0_PERF_WRITE_STALL_SIZE				32


// Register NVDLA_PDP_D_CYA_0
#define NVDLA_PDP_D_CYA_0					32'hb09c
#define NVDLA_PDP_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_PDP_D_CYA_0_CYA_SIZE				32


// Register NVDLA_CDP_RDMA_S_STATUS_0
#define NVDLA_CDP_RDMA_S_STATUS_0					32'hc000
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CDP_RDMA_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CDP_RDMA_S_POINTER_0
#define NVDLA_CDP_RDMA_S_POINTER_0					32'hc004
#define NVDLA_CDP_RDMA_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CDP_RDMA_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CDP_RDMA_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CDP_RDMA_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CDP_RDMA_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CDP_RDMA_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CDP_RDMA_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CDP_RDMA_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CDP_RDMA_D_OP_ENABLE_0
#define NVDLA_CDP_RDMA_D_OP_ENABLE_0					32'hc008
#define NVDLA_CDP_RDMA_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CDP_RDMA_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CDP_RDMA_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CDP_RDMA_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CDP_RDMA_D_DATA_CUBE_WIDTH_0
#define NVDLA_CDP_RDMA_D_DATA_CUBE_WIDTH_0					32'hc00c
#define NVDLA_CDP_RDMA_D_DATA_CUBE_WIDTH_0_WIDTH_RANGE			12:0
#define NVDLA_CDP_RDMA_D_DATA_CUBE_WIDTH_0_WIDTH_SIZE				13


// Register NVDLA_CDP_RDMA_D_DATA_CUBE_HEIGHT_0
#define NVDLA_CDP_RDMA_D_DATA_CUBE_HEIGHT_0					32'hc010
#define NVDLA_CDP_RDMA_D_DATA_CUBE_HEIGHT_0_HEIGHT_RANGE			12:0
#define NVDLA_CDP_RDMA_D_DATA_CUBE_HEIGHT_0_HEIGHT_SIZE				13


// Register NVDLA_CDP_RDMA_D_DATA_CUBE_CHANNEL_0
#define NVDLA_CDP_RDMA_D_DATA_CUBE_CHANNEL_0					32'hc014
#define NVDLA_CDP_RDMA_D_DATA_CUBE_CHANNEL_0_CHANNEL_RANGE			12:0
#define NVDLA_CDP_RDMA_D_DATA_CUBE_CHANNEL_0_CHANNEL_SIZE				13


// Register NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_LOW_0					32'hc018
#define NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_HIGH_0					32'hc01c
#define NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_CDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_CDP_RDMA_D_SRC_LINE_STRIDE_0
#define NVDLA_CDP_RDMA_D_SRC_LINE_STRIDE_0					32'hc020
#define NVDLA_CDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_CDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_CDP_RDMA_D_SRC_SURFACE_STRIDE_0
#define NVDLA_CDP_RDMA_D_SRC_SURFACE_STRIDE_0					32'hc024
#define NVDLA_CDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_CDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_CDP_RDMA_D_SRC_DMA_CFG_0
#define NVDLA_CDP_RDMA_D_SRC_DMA_CFG_0					32'hc028
#define NVDLA_CDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_RANGE			0:0
#define NVDLA_CDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_SIZE				1
#define NVDLA_CDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_CV			1'h0
#define NVDLA_CDP_RDMA_D_SRC_DMA_CFG_0_SRC_RAM_TYPE_MC			1'h1


// Register NVDLA_CDP_RDMA_D_SRC_COMPRESSION_EN_0
#define NVDLA_CDP_RDMA_D_SRC_COMPRESSION_EN_0					32'hc02c
#define NVDLA_CDP_RDMA_D_SRC_COMPRESSION_EN_0_SRC_COMPRESSION_EN_RANGE			0:0
#define NVDLA_CDP_RDMA_D_SRC_COMPRESSION_EN_0_SRC_COMPRESSION_EN_SIZE				1
#define NVDLA_CDP_RDMA_D_SRC_COMPRESSION_EN_0_SRC_COMPRESSION_EN_DISABLE			1'h0
#define NVDLA_CDP_RDMA_D_SRC_COMPRESSION_EN_0_SRC_COMPRESSION_EN_ENABLE			1'h1


// Register NVDLA_CDP_RDMA_D_OPERATION_MODE_0
#define NVDLA_CDP_RDMA_D_OPERATION_MODE_0					32'hc030
#define NVDLA_CDP_RDMA_D_OPERATION_MODE_0_OPERATION_MODE_RANGE			1:0
#define NVDLA_CDP_RDMA_D_OPERATION_MODE_0_OPERATION_MODE_SIZE				2
#define NVDLA_CDP_RDMA_D_OPERATION_MODE_0_OPERATION_MODE_READPHILE			2'h0
#define NVDLA_CDP_RDMA_D_OPERATION_MODE_0_OPERATION_MODE_WRITEPHILE			2'h1
#define NVDLA_CDP_RDMA_D_OPERATION_MODE_0_OPERATION_MODE_ORDINARY			2'h2


// Register NVDLA_CDP_RDMA_D_DATA_FORMAT_0
#define NVDLA_CDP_RDMA_D_DATA_FORMAT_0					32'hc034
#define NVDLA_CDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_RANGE			1:0
#define NVDLA_CDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_SIZE				2
#define NVDLA_CDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_INT8			2'h0
#define NVDLA_CDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_INT16			2'h1
#define NVDLA_CDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_FP16			2'h2


// Register NVDLA_CDP_RDMA_D_PERF_ENABLE_0
#define NVDLA_CDP_RDMA_D_PERF_ENABLE_0					32'hc038
#define NVDLA_CDP_RDMA_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_CDP_RDMA_D_PERF_ENABLE_0_DMA_EN_SIZE				1
#define NVDLA_CDP_RDMA_D_PERF_ENABLE_0_DMA_EN_DISABLE			1'h0
#define NVDLA_CDP_RDMA_D_PERF_ENABLE_0_DMA_EN_ENABLE			1'h1


// Register NVDLA_CDP_RDMA_D_PERF_READ_STALL_0
#define NVDLA_CDP_RDMA_D_PERF_READ_STALL_0					32'hc03c
#define NVDLA_CDP_RDMA_D_PERF_READ_STALL_0_PERF_READ_STALL_RANGE			31:0
#define NVDLA_CDP_RDMA_D_PERF_READ_STALL_0_PERF_READ_STALL_SIZE				32


// Register NVDLA_CDP_RDMA_D_CYA_0
#define NVDLA_CDP_RDMA_D_CYA_0					32'hc040
#define NVDLA_CDP_RDMA_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CDP_RDMA_D_CYA_0_CYA_SIZE				32


// Register NVDLA_CDP_S_STATUS_0
#define NVDLA_CDP_S_STATUS_0					32'hd000
#define NVDLA_CDP_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CDP_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CDP_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CDP_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CDP_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CDP_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CDP_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CDP_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CDP_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CDP_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CDP_S_POINTER_0
#define NVDLA_CDP_S_POINTER_0					32'hd004
#define NVDLA_CDP_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CDP_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CDP_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CDP_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CDP_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CDP_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CDP_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CDP_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CDP_S_LUT_ACCESS_CFG_0
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0					32'hd008
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_ADDR_RANGE			9:0
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_ADDR_SIZE				10
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_RANGE			16:16
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_SIZE				1
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_LE			1'h0
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_LO			1'h1
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_RANGE			17:17
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_SIZE				1
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_READ			1'h0
#define NVDLA_CDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_WRITE			1'h1


// Register NVDLA_CDP_S_LUT_ACCESS_DATA_0
#define NVDLA_CDP_S_LUT_ACCESS_DATA_0					32'hd00c
#define NVDLA_CDP_S_LUT_ACCESS_DATA_0_LUT_DATA_RANGE			15:0
#define NVDLA_CDP_S_LUT_ACCESS_DATA_0_LUT_DATA_SIZE				16


// Register NVDLA_CDP_S_LUT_CFG_0
#define NVDLA_CDP_S_LUT_CFG_0					32'hd010
#define NVDLA_CDP_S_LUT_CFG_0_LUT_LE_FUNCTION_RANGE			0:0
#define NVDLA_CDP_S_LUT_CFG_0_LUT_LE_FUNCTION_SIZE				1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_LE_FUNCTION_EXPONENT			1'h0
#define NVDLA_CDP_S_LUT_CFG_0_LUT_LE_FUNCTION_LINEAR			1'h1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_RANGE			4:4
#define NVDLA_CDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_SIZE				1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_LE			1'h0
#define NVDLA_CDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_LO			1'h1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_RANGE			5:5
#define NVDLA_CDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_SIZE				1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_LE			1'h0
#define NVDLA_CDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_LO			1'h1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_RANGE			6:6
#define NVDLA_CDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_SIZE				1
#define NVDLA_CDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_LE			1'h0
#define NVDLA_CDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_LO			1'h1


// Register NVDLA_CDP_S_LUT_INFO_0
#define NVDLA_CDP_S_LUT_INFO_0					32'hd014
#define NVDLA_CDP_S_LUT_INFO_0_LUT_LE_INDEX_OFFSET_RANGE			7:0
#define NVDLA_CDP_S_LUT_INFO_0_LUT_LE_INDEX_OFFSET_SIZE				8
#define NVDLA_CDP_S_LUT_INFO_0_LUT_LE_INDEX_SELECT_RANGE			15:8
#define NVDLA_CDP_S_LUT_INFO_0_LUT_LE_INDEX_SELECT_SIZE				8
#define NVDLA_CDP_S_LUT_INFO_0_LUT_LO_INDEX_SELECT_RANGE			23:16
#define NVDLA_CDP_S_LUT_INFO_0_LUT_LO_INDEX_SELECT_SIZE				8


// Register NVDLA_CDP_S_LUT_LE_START_LOW_0
#define NVDLA_CDP_S_LUT_LE_START_LOW_0					32'hd018
#define NVDLA_CDP_S_LUT_LE_START_LOW_0_LUT_LE_START_LOW_RANGE			31:0
#define NVDLA_CDP_S_LUT_LE_START_LOW_0_LUT_LE_START_LOW_SIZE				32


// Register NVDLA_CDP_S_LUT_LE_START_HIGH_0
#define NVDLA_CDP_S_LUT_LE_START_HIGH_0					32'hd01c
#define NVDLA_CDP_S_LUT_LE_START_HIGH_0_LUT_LE_START_HIGH_RANGE			5:0
#define NVDLA_CDP_S_LUT_LE_START_HIGH_0_LUT_LE_START_HIGH_SIZE				6


// Register NVDLA_CDP_S_LUT_LE_END_LOW_0
#define NVDLA_CDP_S_LUT_LE_END_LOW_0					32'hd020
#define NVDLA_CDP_S_LUT_LE_END_LOW_0_LUT_LE_END_LOW_RANGE			31:0
#define NVDLA_CDP_S_LUT_LE_END_LOW_0_LUT_LE_END_LOW_SIZE				32


// Register NVDLA_CDP_S_LUT_LE_END_HIGH_0
#define NVDLA_CDP_S_LUT_LE_END_HIGH_0					32'hd024
#define NVDLA_CDP_S_LUT_LE_END_HIGH_0_LUT_LE_END_HIGH_RANGE			5:0
#define NVDLA_CDP_S_LUT_LE_END_HIGH_0_LUT_LE_END_HIGH_SIZE				6


// Register NVDLA_CDP_S_LUT_LO_START_LOW_0
#define NVDLA_CDP_S_LUT_LO_START_LOW_0					32'hd028
#define NVDLA_CDP_S_LUT_LO_START_LOW_0_LUT_LO_START_LOW_RANGE			31:0
#define NVDLA_CDP_S_LUT_LO_START_LOW_0_LUT_LO_START_LOW_SIZE				32


// Register NVDLA_CDP_S_LUT_LO_START_HIGH_0
#define NVDLA_CDP_S_LUT_LO_START_HIGH_0					32'hd02c
#define NVDLA_CDP_S_LUT_LO_START_HIGH_0_LUT_LO_START_HIGH_RANGE			5:0
#define NVDLA_CDP_S_LUT_LO_START_HIGH_0_LUT_LO_START_HIGH_SIZE				6


// Register NVDLA_CDP_S_LUT_LO_END_LOW_0
#define NVDLA_CDP_S_LUT_LO_END_LOW_0					32'hd030
#define NVDLA_CDP_S_LUT_LO_END_LOW_0_LUT_LO_END_LOW_RANGE			31:0
#define NVDLA_CDP_S_LUT_LO_END_LOW_0_LUT_LO_END_LOW_SIZE				32


// Register NVDLA_CDP_S_LUT_LO_END_HIGH_0
#define NVDLA_CDP_S_LUT_LO_END_HIGH_0					32'hd034
#define NVDLA_CDP_S_LUT_LO_END_HIGH_0_LUT_LO_END_HIGH_RANGE			5:0
#define NVDLA_CDP_S_LUT_LO_END_HIGH_0_LUT_LO_END_HIGH_SIZE				6


// Register NVDLA_CDP_S_LUT_LE_SLOPE_SCALE_0
#define NVDLA_CDP_S_LUT_LE_SLOPE_SCALE_0					32'hd038
#define NVDLA_CDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_UFLOW_SCALE_RANGE			15:0
#define NVDLA_CDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_UFLOW_SCALE_SIZE				16
#define NVDLA_CDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_OFLOW_SCALE_RANGE			31:16
#define NVDLA_CDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_OFLOW_SCALE_SIZE				16


// Register NVDLA_CDP_S_LUT_LE_SLOPE_SHIFT_0
#define NVDLA_CDP_S_LUT_LE_SLOPE_SHIFT_0					32'hd03c
#define NVDLA_CDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_UFLOW_SHIFT_RANGE			4:0
#define NVDLA_CDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_UFLOW_SHIFT_SIZE				5
#define NVDLA_CDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_OFLOW_SHIFT_RANGE			9:5
#define NVDLA_CDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_OFLOW_SHIFT_SIZE				5


// Register NVDLA_CDP_S_LUT_LO_SLOPE_SCALE_0
#define NVDLA_CDP_S_LUT_LO_SLOPE_SCALE_0					32'hd040
#define NVDLA_CDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_UFLOW_SCALE_RANGE			15:0
#define NVDLA_CDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_UFLOW_SCALE_SIZE				16
#define NVDLA_CDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_OFLOW_SCALE_RANGE			31:16
#define NVDLA_CDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_OFLOW_SCALE_SIZE				16


// Register NVDLA_CDP_S_LUT_LO_SLOPE_SHIFT_0
#define NVDLA_CDP_S_LUT_LO_SLOPE_SHIFT_0					32'hd044
#define NVDLA_CDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_UFLOW_SHIFT_RANGE			4:0
#define NVDLA_CDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_UFLOW_SHIFT_SIZE				5
#define NVDLA_CDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_OFLOW_SHIFT_RANGE			9:5
#define NVDLA_CDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_OFLOW_SHIFT_SIZE				5


// Register NVDLA_CDP_D_OP_ENABLE_0
#define NVDLA_CDP_D_OP_ENABLE_0					32'hd048
#define NVDLA_CDP_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CDP_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CDP_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CDP_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CDP_D_FUNC_BYPASS_0
#define NVDLA_CDP_D_FUNC_BYPASS_0					32'hd04c
#define NVDLA_CDP_D_FUNC_BYPASS_0_SQSUM_BYPASS_RANGE			0:0
#define NVDLA_CDP_D_FUNC_BYPASS_0_SQSUM_BYPASS_SIZE				1
#define NVDLA_CDP_D_FUNC_BYPASS_0_SQSUM_BYPASS_DISABLE			1'h0
#define NVDLA_CDP_D_FUNC_BYPASS_0_SQSUM_BYPASS_ENABLE			1'h1
#define NVDLA_CDP_D_FUNC_BYPASS_0_MUL_BYPASS_RANGE			1:1
#define NVDLA_CDP_D_FUNC_BYPASS_0_MUL_BYPASS_SIZE				1
#define NVDLA_CDP_D_FUNC_BYPASS_0_MUL_BYPASS_DISABLE			1'h0
#define NVDLA_CDP_D_FUNC_BYPASS_0_MUL_BYPASS_ENABLE			1'h1


// Register NVDLA_CDP_D_DST_BASE_ADDR_LOW_0
#define NVDLA_CDP_D_DST_BASE_ADDR_LOW_0					32'hd050
#define NVDLA_CDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_CDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_CDP_D_DST_BASE_ADDR_HIGH_0
#define NVDLA_CDP_D_DST_BASE_ADDR_HIGH_0					32'hd054
#define NVDLA_CDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_CDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_CDP_D_DST_LINE_STRIDE_0
#define NVDLA_CDP_D_DST_LINE_STRIDE_0					32'hd058
#define NVDLA_CDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_RANGE			31:0
#define NVDLA_CDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_SIZE				32


// Register NVDLA_CDP_D_DST_SURFACE_STRIDE_0
#define NVDLA_CDP_D_DST_SURFACE_STRIDE_0					32'hd05c
#define NVDLA_CDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_CDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_SIZE				32


// Register NVDLA_CDP_D_DST_DMA_CFG_0
#define NVDLA_CDP_D_DST_DMA_CFG_0					32'hd060
#define NVDLA_CDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_RANGE			0:0
#define NVDLA_CDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_SIZE				1
#define NVDLA_CDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_CV			1'h0
#define NVDLA_CDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_MC			1'h1


// Register NVDLA_CDP_D_DST_COMPRESSION_EN_0
#define NVDLA_CDP_D_DST_COMPRESSION_EN_0					32'hd064
#define NVDLA_CDP_D_DST_COMPRESSION_EN_0_DST_COMPRESSION_EN_RANGE			0:0
#define NVDLA_CDP_D_DST_COMPRESSION_EN_0_DST_COMPRESSION_EN_SIZE				1
#define NVDLA_CDP_D_DST_COMPRESSION_EN_0_DST_COMPRESSION_EN_DISABLE			1'h0
#define NVDLA_CDP_D_DST_COMPRESSION_EN_0_DST_COMPRESSION_EN_ENABLE			1'h1


// Register NVDLA_CDP_D_DATA_FORMAT_0
#define NVDLA_CDP_D_DATA_FORMAT_0					32'hd068
#define NVDLA_CDP_D_DATA_FORMAT_0_INPUT_DATA_TYPE_RANGE			1:0
#define NVDLA_CDP_D_DATA_FORMAT_0_INPUT_DATA_TYPE_SIZE				2
#define NVDLA_CDP_D_DATA_FORMAT_0_INPUT_DATA_TYPE_INT8			2'h0
#define NVDLA_CDP_D_DATA_FORMAT_0_INPUT_DATA_TYPE_INT16			2'h1
#define NVDLA_CDP_D_DATA_FORMAT_0_INPUT_DATA_TYPE_FP16			2'h2


// Register NVDLA_CDP_D_NAN_FLUSH_TO_ZERO_0
#define NVDLA_CDP_D_NAN_FLUSH_TO_ZERO_0					32'hd06c
#define NVDLA_CDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_RANGE			0:0
#define NVDLA_CDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_SIZE				1
#define NVDLA_CDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_DISABLE			1'h0
#define NVDLA_CDP_D_NAN_FLUSH_TO_ZERO_0_NAN_TO_ZERO_ENABLE			1'h1


// Register NVDLA_CDP_D_LRN_CFG_0
#define NVDLA_CDP_D_LRN_CFG_0					32'hd070
#define NVDLA_CDP_D_LRN_CFG_0_NORMALZ_LEN_RANGE			1:0
#define NVDLA_CDP_D_LRN_CFG_0_NORMALZ_LEN_SIZE				2
#define NVDLA_CDP_D_LRN_CFG_0_NORMALZ_LEN_LEN3			2'h0
#define NVDLA_CDP_D_LRN_CFG_0_NORMALZ_LEN_LEN5			2'h1
#define NVDLA_CDP_D_LRN_CFG_0_NORMALZ_LEN_LEN7			2'h2
#define NVDLA_CDP_D_LRN_CFG_0_NORMALZ_LEN_LEN9			2'h3


// Register NVDLA_CDP_D_DATIN_OFFSET_0
#define NVDLA_CDP_D_DATIN_OFFSET_0					32'hd074
#define NVDLA_CDP_D_DATIN_OFFSET_0_DATIN_OFFSET_RANGE			15:0
#define NVDLA_CDP_D_DATIN_OFFSET_0_DATIN_OFFSET_SIZE				16


// Register NVDLA_CDP_D_DATIN_SCALE_0
#define NVDLA_CDP_D_DATIN_SCALE_0					32'hd078
#define NVDLA_CDP_D_DATIN_SCALE_0_DATIN_SCALE_RANGE			15:0
#define NVDLA_CDP_D_DATIN_SCALE_0_DATIN_SCALE_SIZE				16


// Register NVDLA_CDP_D_DATIN_SHIFTER_0
#define NVDLA_CDP_D_DATIN_SHIFTER_0					32'hd07c
#define NVDLA_CDP_D_DATIN_SHIFTER_0_DATIN_SHIFTER_RANGE			4:0
#define NVDLA_CDP_D_DATIN_SHIFTER_0_DATIN_SHIFTER_SIZE				5


// Register NVDLA_CDP_D_DATOUT_OFFSET_0
#define NVDLA_CDP_D_DATOUT_OFFSET_0					32'hd080
#define NVDLA_CDP_D_DATOUT_OFFSET_0_DATOUT_OFFSET_RANGE			31:0
#define NVDLA_CDP_D_DATOUT_OFFSET_0_DATOUT_OFFSET_SIZE				32


// Register NVDLA_CDP_D_DATOUT_SCALE_0
#define NVDLA_CDP_D_DATOUT_SCALE_0					32'hd084
#define NVDLA_CDP_D_DATOUT_SCALE_0_DATOUT_SCALE_RANGE			15:0
#define NVDLA_CDP_D_DATOUT_SCALE_0_DATOUT_SCALE_SIZE				16


// Register NVDLA_CDP_D_DATOUT_SHIFTER_0
#define NVDLA_CDP_D_DATOUT_SHIFTER_0					32'hd088
#define NVDLA_CDP_D_DATOUT_SHIFTER_0_DATOUT_SHIFTER_RANGE			5:0
#define NVDLA_CDP_D_DATOUT_SHIFTER_0_DATOUT_SHIFTER_SIZE				6


// Register NVDLA_CDP_D_NAN_INPUT_NUM_0
#define NVDLA_CDP_D_NAN_INPUT_NUM_0					32'hd08c
#define NVDLA_CDP_D_NAN_INPUT_NUM_0_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_CDP_D_NAN_INPUT_NUM_0_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_CDP_D_INF_INPUT_NUM_0
#define NVDLA_CDP_D_INF_INPUT_NUM_0					32'hd090
#define NVDLA_CDP_D_INF_INPUT_NUM_0_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_CDP_D_INF_INPUT_NUM_0_INF_INPUT_NUM_SIZE				32


// Register NVDLA_CDP_D_NAN_OUTPUT_NUM_0
#define NVDLA_CDP_D_NAN_OUTPUT_NUM_0					32'hd094
#define NVDLA_CDP_D_NAN_OUTPUT_NUM_0_NAN_OUTPUT_NUM_RANGE			31:0
#define NVDLA_CDP_D_NAN_OUTPUT_NUM_0_NAN_OUTPUT_NUM_SIZE				32


// Register NVDLA_CDP_D_OUT_SATURATION_0
#define NVDLA_CDP_D_OUT_SATURATION_0					32'hd098
#define NVDLA_CDP_D_OUT_SATURATION_0_OUT_SATURATION_RANGE			31:0
#define NVDLA_CDP_D_OUT_SATURATION_0_OUT_SATURATION_SIZE				32


// Register NVDLA_CDP_D_PERF_ENABLE_0
#define NVDLA_CDP_D_PERF_ENABLE_0					32'hd09c
#define NVDLA_CDP_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_CDP_D_PERF_ENABLE_0_DMA_EN_SIZE				1
#define NVDLA_CDP_D_PERF_ENABLE_0_DMA_EN_DISABLE			1'h0
#define NVDLA_CDP_D_PERF_ENABLE_0_DMA_EN_ENABLE			1'h1
#define NVDLA_CDP_D_PERF_ENABLE_0_LUT_EN_RANGE			1:1
#define NVDLA_CDP_D_PERF_ENABLE_0_LUT_EN_SIZE				1
#define NVDLA_CDP_D_PERF_ENABLE_0_LUT_EN_DISABLE			1'h0
#define NVDLA_CDP_D_PERF_ENABLE_0_LUT_EN_ENABLE			1'h1


// Register NVDLA_CDP_D_PERF_WRITE_STALL_0
#define NVDLA_CDP_D_PERF_WRITE_STALL_0					32'hd0a0
#define NVDLA_CDP_D_PERF_WRITE_STALL_0_PERF_WRITE_STALL_RANGE			31:0
#define NVDLA_CDP_D_PERF_WRITE_STALL_0_PERF_WRITE_STALL_SIZE				32


// Register NVDLA_CDP_D_PERF_LUT_UFLOW_0
#define NVDLA_CDP_D_PERF_LUT_UFLOW_0					32'hd0a4
#define NVDLA_CDP_D_PERF_LUT_UFLOW_0_PERF_LUT_UFLOW_RANGE			31:0
#define NVDLA_CDP_D_PERF_LUT_UFLOW_0_PERF_LUT_UFLOW_SIZE				32


// Register NVDLA_CDP_D_PERF_LUT_OFLOW_0
#define NVDLA_CDP_D_PERF_LUT_OFLOW_0					32'hd0a8
#define NVDLA_CDP_D_PERF_LUT_OFLOW_0_PERF_LUT_OFLOW_RANGE			31:0
#define NVDLA_CDP_D_PERF_LUT_OFLOW_0_PERF_LUT_OFLOW_SIZE				32


// Register NVDLA_CDP_D_PERF_LUT_HYBRID_0
#define NVDLA_CDP_D_PERF_LUT_HYBRID_0					32'hd0ac
#define NVDLA_CDP_D_PERF_LUT_HYBRID_0_PERF_LUT_HYBRID_RANGE			31:0
#define NVDLA_CDP_D_PERF_LUT_HYBRID_0_PERF_LUT_HYBRID_SIZE				32


// Register NVDLA_CDP_D_PERF_LUT_LE_HIT_0
#define NVDLA_CDP_D_PERF_LUT_LE_HIT_0					32'hd0b0
#define NVDLA_CDP_D_PERF_LUT_LE_HIT_0_PERF_LUT_LE_HIT_RANGE			31:0
#define NVDLA_CDP_D_PERF_LUT_LE_HIT_0_PERF_LUT_LE_HIT_SIZE				32


// Register NVDLA_CDP_D_PERF_LUT_LO_HIT_0
#define NVDLA_CDP_D_PERF_LUT_LO_HIT_0					32'hd0b4
#define NVDLA_CDP_D_PERF_LUT_LO_HIT_0_PERF_LUT_LO_HIT_RANGE			31:0
#define NVDLA_CDP_D_PERF_LUT_LO_HIT_0_PERF_LUT_LO_HIT_SIZE				32


// Register NVDLA_CDP_D_CYA_0
#define NVDLA_CDP_D_CYA_0					32'hd0b8
#define NVDLA_CDP_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CDP_D_CYA_0_CYA_SIZE				32


// Register NVDLA_GEC_FEATURE_0
#define NVDLA_GEC_FEATURE_0					32'he000
#define NVDLA_GEC_FEATURE_0_NUM_ERR_SLICES_RANGE			5:0
#define NVDLA_GEC_FEATURE_0_NUM_ERR_SLICES_SIZE				6
#define NVDLA_GEC_FEATURE_0_NUM_ERR_RANGE			31:16
#define NVDLA_GEC_FEATURE_0_NUM_ERR_SIZE				16


// Register NVDLA_GEC_SWRESET_0
#define NVDLA_GEC_SWRESET_0					32'he004
#define NVDLA_GEC_SWRESET_0_SWRST_RANGE			0:0
#define NVDLA_GEC_SWRESET_0_SWRST_SIZE				1


// Register NVDLA_GEC_MISSIONERR_TYPE_0
#define NVDLA_GEC_MISSIONERR_TYPE_0					32'he008
#define NVDLA_GEC_MISSIONERR_TYPE_0_CODE_RANGE			5:0
#define NVDLA_GEC_MISSIONERR_TYPE_0_CODE_SIZE				6


// Register NVDLA_GEC_CURRENT_COUNTER_VALUE_0
#define NVDLA_GEC_CURRENT_COUNTER_VALUE_0					32'he00c
#define NVDLA_GEC_CURRENT_COUNTER_VALUE_0_VALUE_RANGE			8:0
#define NVDLA_GEC_CURRENT_COUNTER_VALUE_0_VALUE_SIZE				9


// Register NVDLA_GEC_MISSIONERR_INDEX_0
#define NVDLA_GEC_MISSIONERR_INDEX_0					32'he014
#define NVDLA_GEC_MISSIONERR_INDEX_0_IDX_RANGE			6:0
#define NVDLA_GEC_MISSIONERR_INDEX_0_IDX_SIZE				7


// Register NVDLA_GEC_CORRECTABLE_THRESHOLD_0
#define NVDLA_GEC_CORRECTABLE_THRESHOLD_0					32'he018
#define NVDLA_GEC_CORRECTABLE_THRESHOLD_0_COUNT_RANGE			7:0
#define NVDLA_GEC_CORRECTABLE_THRESHOLD_0_COUNT_SIZE				8


// Register NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0					32'he01c
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_RANGE			7:0
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_SIZE				8
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_LOCK			8'h0
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_UNLOCK			8'he1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0					32'he030
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0					32'he034
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0					32'he038
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR31_SIZE				1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0					32'he03c
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0					32'he040
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0					32'he044
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0					32'he048
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR31_SIZE				1


// Register NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0					32'he050
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_RELOAD			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0					32'he060
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0					32'he064
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0					32'he068
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR63_SIZE				1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0					32'he06c
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0					32'he070
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0					32'he074
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0					32'he078
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR63_SIZE				1


// Register NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0					32'he080
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_RELOAD			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0					32'he084
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0					32'he090
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0					32'he094
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0					32'he098
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR67_SIZE				1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0					32'he09c
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0					32'he0a0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0					32'he0a4
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0					32'he0a8
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR67_SIZE				1


// Register NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0					32'he0b0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_RELOAD			1'h1


// Register NVDLA_CVIF_CFG_RD_WEIGHT_0_0
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0					32'hf000
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_BDMA_RANGE			7:0
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_BDMA_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_SDP_RANGE			15:8
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_SDP_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_PDP_RANGE			23:16
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_PDP_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_CDP_RANGE			31:24
#define NVDLA_CVIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_CDP_SIZE				8


// Register NVDLA_CVIF_CFG_RD_WEIGHT_1_0
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0					32'hf004
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_B_RANGE			7:0
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_B_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_N_RANGE			15:8
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_N_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_E_RANGE			23:16
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_E_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_CDMA_DAT_RANGE			31:24
#define NVDLA_CVIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_CDMA_DAT_SIZE				8


// Register NVDLA_CVIF_CFG_RD_WEIGHT_2_0
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0					32'hf008
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_CDMA_WT_RANGE			7:0
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_CDMA_WT_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RBK_RANGE			15:8
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RBK_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_1_RANGE			23:16
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_1_SIZE				8
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_0_RANGE			31:24
#define NVDLA_CVIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_0_SIZE				8


// Register NVDLA_CVIF_CFG_WR_WEIGHT_0_0
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0					32'hf00c
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_BDMA_RANGE			7:0
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_BDMA_SIZE				8
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_SDP_RANGE			15:8
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_SDP_SIZE				8
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_PDP_RANGE			23:16
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_PDP_SIZE				8
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_CDP_RANGE			31:24
#define NVDLA_CVIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_CDP_SIZE				8


// Register NVDLA_CVIF_CFG_WR_WEIGHT_1_0
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0					32'hf010
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RBK_RANGE			7:0
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RBK_SIZE				8
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_2_RANGE			15:8
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_2_SIZE				8
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_1_RANGE			23:16
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_1_SIZE				8
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_0_RANGE			31:24
#define NVDLA_CVIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_0_SIZE				8


// Register NVDLA_CVIF_CFG_OUTSTANDING_CNT_0
#define NVDLA_CVIF_CFG_OUTSTANDING_CNT_0					32'hf014
#define NVDLA_CVIF_CFG_OUTSTANDING_CNT_0_RD_OS_CNT_RANGE			7:0
#define NVDLA_CVIF_CFG_OUTSTANDING_CNT_0_RD_OS_CNT_SIZE				8
#define NVDLA_CVIF_CFG_OUTSTANDING_CNT_0_WR_OS_CNT_RANGE			15:8
#define NVDLA_CVIF_CFG_OUTSTANDING_CNT_0_WR_OS_CNT_SIZE				8


// Register NVDLA_CVIF_STATUS_0
#define NVDLA_CVIF_STATUS_0					32'hf018
#define NVDLA_CVIF_STATUS_0_IDLE_RANGE			8:8
#define NVDLA_CVIF_STATUS_0_IDLE_SIZE				1
#define NVDLA_CVIF_STATUS_0_IDLE_NO			1'h0
#define NVDLA_CVIF_STATUS_0_IDLE_YES			1'h1


// Register NVDLA_BDMA_CFG_SRC_ADDR_LOW_0
#define NVDLA_BDMA_CFG_SRC_ADDR_LOW_0					32'h10000
#define NVDLA_BDMA_CFG_SRC_ADDR_LOW_0_V32_RANGE			31:5
#define NVDLA_BDMA_CFG_SRC_ADDR_LOW_0_V32_SIZE				27


// Register NVDLA_BDMA_CFG_SRC_ADDR_HIGH_0
#define NVDLA_BDMA_CFG_SRC_ADDR_HIGH_0					32'h10004
#define NVDLA_BDMA_CFG_SRC_ADDR_HIGH_0_V8_RANGE			31:0
#define NVDLA_BDMA_CFG_SRC_ADDR_HIGH_0_V8_SIZE				32


// Register NVDLA_BDMA_CFG_DST_ADDR_LOW_0
#define NVDLA_BDMA_CFG_DST_ADDR_LOW_0					32'h10008
#define NVDLA_BDMA_CFG_DST_ADDR_LOW_0_V32_RANGE			31:5
#define NVDLA_BDMA_CFG_DST_ADDR_LOW_0_V32_SIZE				27


// Register NVDLA_BDMA_CFG_DST_ADDR_HIGH_0
#define NVDLA_BDMA_CFG_DST_ADDR_HIGH_0					32'h1000c
#define NVDLA_BDMA_CFG_DST_ADDR_HIGH_0_V8_RANGE			31:0
#define NVDLA_BDMA_CFG_DST_ADDR_HIGH_0_V8_SIZE				32


// Register NVDLA_BDMA_CFG_LINE_0
#define NVDLA_BDMA_CFG_LINE_0					32'h10010
#define NVDLA_BDMA_CFG_LINE_0_SIZE_RANGE			12:0
#define NVDLA_BDMA_CFG_LINE_0_SIZE_SIZE				13


// Register NVDLA_BDMA_CFG_CMD_0
#define NVDLA_BDMA_CFG_CMD_0					32'h10014
#define NVDLA_BDMA_CFG_CMD_0_SRC_RAM_TYPE_RANGE			0:0
#define NVDLA_BDMA_CFG_CMD_0_SRC_RAM_TYPE_SIZE				1
#define NVDLA_BDMA_CFG_CMD_0_SRC_RAM_TYPE_CVSRAM			1'h0
#define NVDLA_BDMA_CFG_CMD_0_SRC_RAM_TYPE_MC			1'h1
#define NVDLA_BDMA_CFG_CMD_0_DST_RAM_TYPE_RANGE			1:1
#define NVDLA_BDMA_CFG_CMD_0_DST_RAM_TYPE_SIZE				1
#define NVDLA_BDMA_CFG_CMD_0_DST_RAM_TYPE_CVSRAM			1'h0
#define NVDLA_BDMA_CFG_CMD_0_DST_RAM_TYPE_MC			1'h1


// Register NVDLA_BDMA_CFG_LINE_REPEAT_0
#define NVDLA_BDMA_CFG_LINE_REPEAT_0					32'h10018
#define NVDLA_BDMA_CFG_LINE_REPEAT_0_NUMBER_RANGE			23:0
#define NVDLA_BDMA_CFG_LINE_REPEAT_0_NUMBER_SIZE				24


// Register NVDLA_BDMA_CFG_SRC_LINE_0
#define NVDLA_BDMA_CFG_SRC_LINE_0					32'h1001c
#define NVDLA_BDMA_CFG_SRC_LINE_0_STRIDE_RANGE			31:5
#define NVDLA_BDMA_CFG_SRC_LINE_0_STRIDE_SIZE				27


// Register NVDLA_BDMA_CFG_DST_LINE_0
#define NVDLA_BDMA_CFG_DST_LINE_0					32'h10020
#define NVDLA_BDMA_CFG_DST_LINE_0_STRIDE_RANGE			31:5
#define NVDLA_BDMA_CFG_DST_LINE_0_STRIDE_SIZE				27


// Register NVDLA_BDMA_CFG_SURF_REPEAT_0
#define NVDLA_BDMA_CFG_SURF_REPEAT_0					32'h10024
#define NVDLA_BDMA_CFG_SURF_REPEAT_0_NUMBER_RANGE			23:0
#define NVDLA_BDMA_CFG_SURF_REPEAT_0_NUMBER_SIZE				24


// Register NVDLA_BDMA_CFG_SRC_SURF_0
#define NVDLA_BDMA_CFG_SRC_SURF_0					32'h10028
#define NVDLA_BDMA_CFG_SRC_SURF_0_STRIDE_RANGE			31:5
#define NVDLA_BDMA_CFG_SRC_SURF_0_STRIDE_SIZE				27


// Register NVDLA_BDMA_CFG_DST_SURF_0
#define NVDLA_BDMA_CFG_DST_SURF_0					32'h1002c
#define NVDLA_BDMA_CFG_DST_SURF_0_STRIDE_RANGE			31:5
#define NVDLA_BDMA_CFG_DST_SURF_0_STRIDE_SIZE				27


// Register NVDLA_BDMA_CFG_OP_0
#define NVDLA_BDMA_CFG_OP_0					32'h10030
#define NVDLA_BDMA_CFG_OP_0_EN_RANGE			0:0
#define NVDLA_BDMA_CFG_OP_0_EN_SIZE				1
#define NVDLA_BDMA_CFG_OP_0_EN_DISABLE			1'h0
#define NVDLA_BDMA_CFG_OP_0_EN_ENABLE			1'h1


// Register NVDLA_BDMA_CFG_LAUNCH0_0
#define NVDLA_BDMA_CFG_LAUNCH0_0					32'h10034
#define NVDLA_BDMA_CFG_LAUNCH0_0_GRP0_LAUNCH_RANGE			0:0
#define NVDLA_BDMA_CFG_LAUNCH0_0_GRP0_LAUNCH_SIZE				1
#define NVDLA_BDMA_CFG_LAUNCH0_0_GRP0_LAUNCH_NO			1'h0
#define NVDLA_BDMA_CFG_LAUNCH0_0_GRP0_LAUNCH_YES			1'h1


// Register NVDLA_BDMA_CFG_LAUNCH1_0
#define NVDLA_BDMA_CFG_LAUNCH1_0					32'h10038
#define NVDLA_BDMA_CFG_LAUNCH1_0_GRP1_LAUNCH_RANGE			0:0
#define NVDLA_BDMA_CFG_LAUNCH1_0_GRP1_LAUNCH_SIZE				1
#define NVDLA_BDMA_CFG_LAUNCH1_0_GRP1_LAUNCH_NO			1'h0
#define NVDLA_BDMA_CFG_LAUNCH1_0_GRP1_LAUNCH_YES			1'h1


// Register NVDLA_BDMA_CFG_STATUS_0
#define NVDLA_BDMA_CFG_STATUS_0					32'h1003c
#define NVDLA_BDMA_CFG_STATUS_0_STALL_COUNT_EN_RANGE			0:0
#define NVDLA_BDMA_CFG_STATUS_0_STALL_COUNT_EN_SIZE				1
#define NVDLA_BDMA_CFG_STATUS_0_STALL_COUNT_EN_NO			1'h0
#define NVDLA_BDMA_CFG_STATUS_0_STALL_COUNT_EN_YES			1'h1


// Register NVDLA_BDMA_STATUS_0
#define NVDLA_BDMA_STATUS_0					32'h10040
#define NVDLA_BDMA_STATUS_0_FREE_SLOT_RANGE			7:0
#define NVDLA_BDMA_STATUS_0_FREE_SLOT_SIZE				8
#define NVDLA_BDMA_STATUS_0_IDLE_RANGE			8:8
#define NVDLA_BDMA_STATUS_0_IDLE_SIZE				1
#define NVDLA_BDMA_STATUS_0_IDLE_NO			1'h0
#define NVDLA_BDMA_STATUS_0_IDLE_YES			1'h1
#define NVDLA_BDMA_STATUS_0_GRP0_BUSY_RANGE			9:9
#define NVDLA_BDMA_STATUS_0_GRP0_BUSY_SIZE				1
#define NVDLA_BDMA_STATUS_0_GRP0_BUSY_NO			1'h0
#define NVDLA_BDMA_STATUS_0_GRP0_BUSY_YES			1'h1
#define NVDLA_BDMA_STATUS_0_GRP1_BUSY_RANGE			10:10
#define NVDLA_BDMA_STATUS_0_GRP1_BUSY_SIZE				1
#define NVDLA_BDMA_STATUS_0_GRP1_BUSY_NO			1'h0
#define NVDLA_BDMA_STATUS_0_GRP1_BUSY_YES			1'h1


// Register NVDLA_BDMA_STATUS_GRP0_READ_STALL_0
#define NVDLA_BDMA_STATUS_GRP0_READ_STALL_0					32'h10044
#define NVDLA_BDMA_STATUS_GRP0_READ_STALL_0_COUNT_RANGE			31:0
#define NVDLA_BDMA_STATUS_GRP0_READ_STALL_0_COUNT_SIZE				32


// Register NVDLA_BDMA_STATUS_GRP0_WRITE_STALL_0
#define NVDLA_BDMA_STATUS_GRP0_WRITE_STALL_0					32'h10048
#define NVDLA_BDMA_STATUS_GRP0_WRITE_STALL_0_COUNT_RANGE			31:0
#define NVDLA_BDMA_STATUS_GRP0_WRITE_STALL_0_COUNT_SIZE				32


// Register NVDLA_BDMA_STATUS_GRP1_READ_STALL_0
#define NVDLA_BDMA_STATUS_GRP1_READ_STALL_0					32'h1004c
#define NVDLA_BDMA_STATUS_GRP1_READ_STALL_0_COUNT_RANGE			31:0
#define NVDLA_BDMA_STATUS_GRP1_READ_STALL_0_COUNT_SIZE				32


// Register NVDLA_BDMA_STATUS_GRP1_WRITE_STALL_0
#define NVDLA_BDMA_STATUS_GRP1_WRITE_STALL_0					32'h10050
#define NVDLA_BDMA_STATUS_GRP1_WRITE_STALL_0_COUNT_RANGE			31:0
#define NVDLA_BDMA_STATUS_GRP1_WRITE_STALL_0_COUNT_SIZE				32


// Register NVDLA_RBK_S_STATUS_0
#define NVDLA_RBK_S_STATUS_0					32'h11000
#define NVDLA_RBK_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_RBK_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_RBK_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_RBK_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_RBK_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_RBK_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_RBK_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_RBK_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_RBK_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_RBK_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_RBK_S_POINTER_0
#define NVDLA_RBK_S_POINTER_0					32'h11004
#define NVDLA_RBK_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_RBK_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_RBK_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_RBK_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_RBK_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_RBK_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_RBK_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_RBK_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_RBK_D_OP_ENABLE_0
#define NVDLA_RBK_D_OP_ENABLE_0					32'h11008
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_RBK_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_RBK_D_MISC_CFG_0
#define NVDLA_RBK_D_MISC_CFG_0					32'h1100c
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_RANGE			1:0
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_SIZE				2
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_CONTRACT			2'h0
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_SPLIT			2'h1
#define NVDLA_RBK_D_MISC_CFG_0_RUBIK_MODE_MERGE			2'h2
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_RANGE			9:8
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_RBK_D_MISC_CFG_0_IN_PRECISION_FP16			2'h2


// Register NVDLA_RBK_D_DAIN_RAM_TYPE_0
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0					32'h11010
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_RANGE			0:0
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_SIZE				1
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_CVIF			1'h0
#define NVDLA_RBK_D_DAIN_RAM_TYPE_0_DATAIN_RAM_TYPE_MCIF			1'h1


// Register NVDLA_RBK_D_DATAIN_SIZE_0_0
#define NVDLA_RBK_D_DATAIN_SIZE_0_0					32'h11014
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_WIDTH_RANGE			12:0
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_WIDTH_SIZE				13
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_HEIGHT_RANGE			28:16
#define NVDLA_RBK_D_DATAIN_SIZE_0_0_DATAIN_HEIGHT_SIZE				13


// Register NVDLA_RBK_D_DATAIN_SIZE_1_0
#define NVDLA_RBK_D_DATAIN_SIZE_1_0					32'h11018
#define NVDLA_RBK_D_DATAIN_SIZE_1_0_DATAIN_CHANNEL_RANGE			12:0
#define NVDLA_RBK_D_DATAIN_SIZE_1_0_DATAIN_CHANNEL_SIZE				13


// Register NVDLA_RBK_D_DAIN_ADDR_HIGH_0
#define NVDLA_RBK_D_DAIN_ADDR_HIGH_0					32'h1101c
#define NVDLA_RBK_D_DAIN_ADDR_HIGH_0_DAIN_ADDR_HIGH_RANGE			31:0
#define NVDLA_RBK_D_DAIN_ADDR_HIGH_0_DAIN_ADDR_HIGH_SIZE				32


// Register NVDLA_RBK_D_DAIN_ADDR_LOW_0
#define NVDLA_RBK_D_DAIN_ADDR_LOW_0					32'h11020
#define NVDLA_RBK_D_DAIN_ADDR_LOW_0_DAIN_ADDR_LOW_RANGE			31:5
#define NVDLA_RBK_D_DAIN_ADDR_LOW_0_DAIN_ADDR_LOW_SIZE				27


// Register NVDLA_RBK_D_DAIN_LINE_STRIDE_0
#define NVDLA_RBK_D_DAIN_LINE_STRIDE_0					32'h11024
#define NVDLA_RBK_D_DAIN_LINE_STRIDE_0_DAIN_LINE_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAIN_LINE_STRIDE_0_DAIN_LINE_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAIN_SURF_STRIDE_0
#define NVDLA_RBK_D_DAIN_SURF_STRIDE_0					32'h11028
#define NVDLA_RBK_D_DAIN_SURF_STRIDE_0_DAIN_SURF_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAIN_SURF_STRIDE_0_DAIN_SURF_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0
#define NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0					32'h1102c
#define NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0_DAIN_PLANAR_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAIN_PLANAR_STRIDE_0_DAIN_PLANAR_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAOUT_RAM_TYPE_0
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0					32'h11030
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_RANGE			0:0
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_SIZE				1
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_CVIF			1'h0
#define NVDLA_RBK_D_DAOUT_RAM_TYPE_0_DATAOUT_RAM_TYPE_MCIF			1'h1


// Register NVDLA_RBK_D_DATAOUT_SIZE_1_0
#define NVDLA_RBK_D_DATAOUT_SIZE_1_0					32'h11034
#define NVDLA_RBK_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_RANGE			12:0
#define NVDLA_RBK_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_SIZE				13


// Register NVDLA_RBK_D_DAOUT_ADDR_HIGH_0
#define NVDLA_RBK_D_DAOUT_ADDR_HIGH_0					32'h11038
#define NVDLA_RBK_D_DAOUT_ADDR_HIGH_0_DAOUT_ADDR_HIGH_RANGE			31:0
#define NVDLA_RBK_D_DAOUT_ADDR_HIGH_0_DAOUT_ADDR_HIGH_SIZE				32


// Register NVDLA_RBK_D_DAOUT_ADDR_LOW_0
#define NVDLA_RBK_D_DAOUT_ADDR_LOW_0					32'h1103c
#define NVDLA_RBK_D_DAOUT_ADDR_LOW_0_DAOUT_ADDR_LOW_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_ADDR_LOW_0_DAOUT_ADDR_LOW_SIZE				27


// Register NVDLA_RBK_D_DAOUT_LINE_STRIDE_0
#define NVDLA_RBK_D_DAOUT_LINE_STRIDE_0					32'h11040
#define NVDLA_RBK_D_DAOUT_LINE_STRIDE_0_DAOUT_LINE_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_LINE_STRIDE_0_DAOUT_LINE_STRIDE_SIZE				27


// Register NVDLA_RBK_D_CONTRACT_STRIDE_0_0
#define NVDLA_RBK_D_CONTRACT_STRIDE_0_0					32'h11044
#define NVDLA_RBK_D_CONTRACT_STRIDE_0_0_CONTRACT_STRIDE_0_RANGE			31:5
#define NVDLA_RBK_D_CONTRACT_STRIDE_0_0_CONTRACT_STRIDE_0_SIZE				27


// Register NVDLA_RBK_D_CONTRACT_STRIDE_1_0
#define NVDLA_RBK_D_CONTRACT_STRIDE_1_0					32'h11048
#define NVDLA_RBK_D_CONTRACT_STRIDE_1_0_CONTRACT_STRIDE_1_RANGE			31:5
#define NVDLA_RBK_D_CONTRACT_STRIDE_1_0_CONTRACT_STRIDE_1_SIZE				27


// Register NVDLA_RBK_D_DAOUT_SURF_STRIDE_0
#define NVDLA_RBK_D_DAOUT_SURF_STRIDE_0					32'h1104c
#define NVDLA_RBK_D_DAOUT_SURF_STRIDE_0_DAOUT_SURF_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_SURF_STRIDE_0_DAOUT_SURF_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0
#define NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0					32'h11050
#define NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0_DAOUT_PLANAR_STRIDE_RANGE			31:5
#define NVDLA_RBK_D_DAOUT_PLANAR_STRIDE_0_DAOUT_PLANAR_STRIDE_SIZE				27


// Register NVDLA_RBK_D_DECONV_STRIDE_0
#define NVDLA_RBK_D_DECONV_STRIDE_0					32'h11054
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_X_STRIDE_RANGE			4:0
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_X_STRIDE_SIZE				5
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_Y_STRIDE_RANGE			20:16
#define NVDLA_RBK_D_DECONV_STRIDE_0_DECONV_Y_STRIDE_SIZE				5


// Register NVDLA_RBK_D_PERF_ENABLE_0
#define NVDLA_RBK_D_PERF_ENABLE_0					32'h11058
#define NVDLA_RBK_D_PERF_ENABLE_0_PERF_EN_RANGE			0:0
#define NVDLA_RBK_D_PERF_ENABLE_0_PERF_EN_SIZE				1


// Register NVDLA_RBK_D_PERF_READ_STALL_0
#define NVDLA_RBK_D_PERF_READ_STALL_0					32'h1105c
#define NVDLA_RBK_D_PERF_READ_STALL_0_RD_STALL_CNT_RANGE			31:0
#define NVDLA_RBK_D_PERF_READ_STALL_0_RD_STALL_CNT_SIZE				32


// Register NVDLA_RBK_D_PERF_WRITE_STALL_0
#define NVDLA_RBK_D_PERF_WRITE_STALL_0					32'h11060
#define NVDLA_RBK_D_PERF_WRITE_STALL_0_WR_STALL_CNT_RANGE			31:0
#define NVDLA_RBK_D_PERF_WRITE_STALL_0_WR_STALL_CNT_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_CFGROM	32'h0
#define BASE_ADDRESS_NVDLA_GLB	32'h1000
#define BASE_ADDRESS_NVDLA_MCIF	32'h2000
#define BASE_ADDRESS_NVDLA_CDMA	32'h3000
#define BASE_ADDRESS_NVDLA_CSC	32'h4000
#define BASE_ADDRESS_NVDLA_CMAC_A	32'h5000
#define BASE_ADDRESS_NVDLA_CMAC_B	32'h6000
#define BASE_ADDRESS_NVDLA_CACC	32'h7000
#define BASE_ADDRESS_NVDLA_SDP_RDMA	32'h8000
#define BASE_ADDRESS_NVDLA_SDP	32'h9000
#define BASE_ADDRESS_NVDLA_PDP_RDMA	32'ha000
#define BASE_ADDRESS_NVDLA_PDP	32'hb000
#define BASE_ADDRESS_NVDLA_CDP_RDMA	32'hc000
#define BASE_ADDRESS_NVDLA_CDP	32'hd000
#define BASE_ADDRESS_NVDLA_GEC	32'he000
#define BASE_ADDRESS_NVDLA_CVIF	32'hf000
#define BASE_ADDRESS_NVDLA_BDMA	32'h10000
#define BASE_ADDRESS_NVDLA_RBK	32'h11000
