`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MB5N9i8hpnFFDATRaYiC+bZ1XXWlwTdBztDvO8vzpU0tEe1TJe+yh26Rv1EfxYIRN0yyz+knUAwI
sf6Z5x/qXw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nfu3ZpCT98Tv0VxTayspTywP22MqwBSSpgYjuleh2cCZtHJFOgjEKu4jM/uDRz8sbyJ4R3FkS2Vx
qsVQAYsplWo0l6wI/XNAwxN7iHoPXprN/N37aGGUJ80TcxP69mCcwoithMacWAmQHUvTvxONS2iO
yKnXxyBc20hfmkgis/8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jZS0Sg6Iztp4XA/jmLpAvkehOZdjieHl4YtcGfZstPyKmfJvo+GifvqzKY/B11D8M4HNZxH3BO69
G2mHkIB9cvDAH87dOQGv1bcMsBi98QDVy8LYKXt3Rmfu0jtbog1RO8UctUYYuqSeh4UoZIb4aqEf
K3ZxsXvbYe5Lmye+5gQKLCAr/Fz8DodGVhsp7pD94MCqIn2IFIxk4cDngLOOuG24zH2uWUEXbRF+
jqMiwRCpHXzNdxbD3Xt76MIITAQZf7b90MtK6RJOf747rOqvQ0BRarNdjibiXrNTEb+LDP/MVcWq
EZOS3k4WoKrwxT+mRT3jNQHjOGdPHdv+30OX9g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vqo1f1C99iMrWKdw+RduCyDS1cCCq9ezmSOrk/2lIw8ZJ0gr2LrtKNKH4dyjvOQolDBQ1EVxuzkk
xmvfkOOIBi9JdmNqhQALGWloB07N/IJdMdvv76U9EjLLzdmY541XyQ8MURpIS9d9rz6L+K6aclFa
dXENCepih6i+kx7wKM97pXzwbpDK+KX+Ykc4gyZQPEI4RxfFpp54Xh+Oo0hLhd/aUKWgnoSIMLwp
XNStqnyweDmEKpaN7Lho4D33O3MrS4VLklK3vXkmQ2k1PNAY8vRTb+Hz1M/M9iYBrbYUieP9wYdJ
SzAg0Ifn/ws16ZVZfU4IJscAaPY5YSn+wzmN0A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GsBKnSG8T9ZDD7l8k1MMkmNRtyFVDJRW3f31lhoZf/Y5XUDODhZ9pCskXZgdU++mAIRDpK2sIx2/
cXnwqifBbijmgHxErTD5WxCRkKGwYsDRXGYD5UacMoDM7lQmyc+ezcQjiVJNwN/lSOiFItznNkWQ
BMOO/2NwzS3mN1VgMbQdBHJxjxSARHNV/69JnUC8/lRbl83oJ3Ht+/KTzZ4qr7RfhE6uz+mtK1A3
0KLeh3uD2p6rf+VRZAA1dy4o23FdoA8k9mkcdnhIHYfXRRcMxVkbXo0mByYk5NvRUbDanOAJ9kOD
bZ/t/KLmZH77CcP7M5AbY7SBLyTJyrJaQAgIvA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KQJNaMLE4WXIKyN7P/9TNSZx0n3pcRzJsgnstM1oCTb58/V3PdsptAGbFAK+YKIo0gRaG+Mjj764
6TY5IjZtKoeMNbhE8kplDsv/hjFxmQXCmTwbk1yrTLV6tKr/VuXnJQIvSBrfVVJwJ2MjjVgifBu7
yWyUyKxF/xQ42neMUls=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bS7Nbjm49uf44kPEEORdhBjYLbD56K4GTmDRNlhmMdqcSWTk+dMHIxXTwIKiWj3THN732d0HAK4Q
slXhzt965qBVm6XrnxOv4+hFHhjTFfSCBAKf0oZLkW6lPfBz9ceDfA4u15UMglq6ABW8hVO4c8O+
BYAgAKyGafXIo++6D+4egK4dhsfcVWR/v30z+fx+pWPCHGmZKgHZtqDwoRAR9LGh+6pZvdDPbfkp
7faz6ouPBlp3VyFdZ8cwMcujgazd/4MuFtQcyKDzHk0eqrtNpAnr98w1EuM+Ih+6OptW6Iimbu1j
Wz+WpN+F4IUGeyfk6cDn9VEoFkZ+Hbcmv2qGBA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wTfHmVZg9zMaxVvmg6iebdpnTvxKxA3BKnDjDkPoIML9i4glT5T7B8DyEX4E860gxs9gIxvBtIfv
NOlqrnPszMjWmsjm+5ZklupSvjfDTuOAgAWPDkGDzdDnKVrBwkG6qU4O5NS6iODJfcd5upOKTSKG
kYQUqSbcu/MoQsjxG/bLx5PuCOUZ9Ob9r0QYgtP7wxlgOB1dgQyV67/7v6K+sPymajAsPMZOCNtp
0pgxkv+4syAlEnZIKTEHAmThwrY76BAOV2F4H6mf2XYImPumULVIWJaDQdRxsqDQq1Qcm2UpLifo
OCkRY7yE1O0CA/YAsWk2iLUR8nYT4JOqS7FnCA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55776)
`protect data_block
0WVUNBbYhJC+vGgsjZ2lgqh118bS1mYb6mCxclB7zyCfmUyzazZQFnUCKofdbFn6t4X5vB5VshFp
B8Hu5akqRPfhw15GQJtfuiycI6mf2vq7+fhkegoVrBVr6mf68siEPA1zjVxg7mkLA6DtaU4EqGTo
aK5jZZTzwq58MSFRfHfi303g7W0CD3sKmZUiqyGCENeWJtp3/y5/n4SlAr2BCIQ+8prm4Z0yY8Bv
PvcAAT2Z+hpZLGl8hstnZ5MmtFfKVEWY+QvuL5H2WlsNUsTXp17T3+yhVIth2eRyrJZXSGcDjb0e
uox4iXXJDgFnNVmJxC8iZ2CRfdMhrsAapiJP7YZYnmZxEf4qotVRbrw5pkm3cnMJLP7hWg/+DrFZ
LYLCEysnoXq82ME018nOKSvM8FH/+LA6pWc4UdfYx3X66+s9/uYfD6LNOBkfSJKjde6SGYLApDA3
tT1VK5SPQiTiDHKblTbuLmziyUN96t1YvUjntQP5bxRyuRkJQGvqWqdQQ7+NuZiR9JAT7Vat2cF3
SR6iGZQMm1EXMxBgJQZNeZi1xpF9gH7VvGtvr4dtH2VSPgIs0WMhLfi8Qi53LDp72JuZ1p/YOb3H
9GRJtnFjRMvpqU9Tz5Gpxc8MRyrSY2UAPJwvdl7a8jisdMRWbbfDt0w24W9GWS30cFO6Fs9pcJ20
C9q36xcYm+7NbhbdCnNQ5trTNvy2wPf98MAF/vzyNrKOH3YcMSBGfYOETiWP8ZIC8CKpRGInt769
7stl23TmnpInycKYGXus/9UM1/hul+4tAombEThOPAiohO6FSe0OkMwNm+Ehy+wsPZct1cIQsAaw
lnZxwgqP4CIxXLzHENi3YMn6Ls7yk26QxJtCJUNSSv0+vJv4PACaXjFugPIE9bKz1AjSVr6NB7UI
iNCZCiGjKY8yO0HxFUXVYD/vhTVSOSp+3yNl8FXSlgpvQrnP5iT/ZhFJ99U5zk2U8M/Wl/t7XUlO
+x9L0wcMTFqRrtsSuhID4HbkxzBtvWoXbfxxZNeklU9PhrSKN3eoZtZ+cFBXuKSPAI1t9htNUNDZ
/PqMRZwAA36LXRbTDnCQXEsu5bmB5z3wRRRuPAyXmQdxWB5Z9fzxbuOcXph+UYWbIqYgG6zJw60c
O90DBKyC5Jk+E5PG2zBmS+l9+tNWXkY5UwJ7T+QsvKFcabGAPh6VhdIXkm7107k/z2BH5BhTWqoa
r6HAtCYjIoGlQvAnN711OIGNQpYmBqHkKSDyQJKULSQHyaPeiaLFC49oi3kSDE/J7GkssifzGoP8
sKycfSAlmFJ3xtjXbaf5QJUh3xW70A3wkSRxtUq1MXzz9ED5inre9YhrGJoOh2dophhUS+u6K8Y7
N59/Oobevhv7W9ugHnkRyR0fEj1VUgshUSGWT/wHzz+HacvSYHBPOaPmVYFb1dZg+slAfdXTlorw
A0/YXynQqy9se8GwlOol/nDr90cSHOMtZpY8BJpylOUVTivmEJpzadnm3abiFVhNrRvc1riQbZV8
6ffJzLhdpNmZchIKo4lDV7GSmnKZtf7K2H1Bj0VIK/naB9GxuWLJNvhe1QAI/DWaDDvTD3D74fZC
SYXF7sY44jcRUE9d4EB77q8/sAoJ5UjP0mQD99I9tmN2ogj2E5ITKciBa25rpIqoIl6Xr6W2zAgF
YcCwpbHy5/1D5hRWES2S7qKTkl9JF72SqvwajfnDNEp0Hw24Fqu7WpG707WiKNtQUqq6Jv+T9gtk
EKG2yuWtyuMC8VuI6KnUxUtIyByDGp+Qmqs8ZkecW5W4ckb14qQ9MNho+mmASHnSIvvENVowaxXm
+k+uHDlbKJaX5pFnPJPsQeUNfuLGsl2CzVh8yGamKajXurnRkpf/S7rrfTQo+pghyvvQRb8KbVcV
deimQckJE4cdez35aEt4vqXJ28QKgP6800jJr9in0Osdxsf1Ez5WFqfu10XKmpx4WMXF6eDq1+bT
ysA3PhPb6pa/vqEpY2OBlP2nVzhaIfHLtJQAQHKnnpJUWYtRSKqeNinPnVtT1V8jKI/Gt5ghy0XP
AViEt+8H/ILj+PNXzte6L4EzPrk2QI3QsHqzdCZN+cPgTprwibADHK6h9kToUcqwbl7VvE0hFLvd
57EEEcu8n/lTE3C+loZwcfbUCSvic1jDlexeMpTOaxFAiNleEQZ4khx7vzFt5tX75a1rqw3CXkXR
fywFmXQxW+fq628pL8SYqS3/bCIPl0STWD6hmmiZgnEeVPDRb7epmsOMsQOAAYZ2vp6xrXbPk9UH
MHtVGdmfAcZrR0iZrYoNDTfFOQ1oTZPo5z4IxdCylnzAgmnZilJkEJ5YLKZ51A7/Mm3U++McquV4
PWDq3Sjig2q8Q4M/qFGxIvSXN4rHBUvVbbtuObXBodz6s2kLBzlrT7c5I94JoKs9LQOtIk2Qa+v5
9UtNR7HfiudQiI7j5d37FRuWtkOMH1SmabeMvcRTv8ua5oKEZFm+ZXPO84E10HoStBY7pVhuqQYY
Ucqg8mTOmO4IiM3jL0OOuvPf/l8o5+b8DE3vjrmDlyD9w1XEETcMoxjbjWC2yq2x8awEW/BkA1Xi
dZn7azC/VpI06wBL4KE8bjYSkkyAqdN/1ya1BJmaxTqcPGDxm7lg4Vuott1fex0xl+oUftDlPoOR
01a4vCkc6BJY35GIg+pHiWCEFJFStsBYtd+2ZML0oiphoHQQhluxGGkUPbnirEuV1lemzsXHsHeN
3n2fOHqk1+5i71xxEMSiQxYHMG2HnANhaQK27L0sv1kQf0tKquS/sk4Q/xNt1Yit2ze1TAlRA9/2
IRHVE6ucZX9N9S4QVmDiD8+fiJI9BlvnBNxPDweCUvRjloGyLBM5WFuyL1kQPHsnRXupkKgiQVjB
Z2BKSjHv9oC3+Rjh/lUSHyNmh06wB7aUpPU6TpNP2CR/ACaubdasVJLqE7X6vQK/covMfxcHLZig
2EzviHWETy49WpfYjzrVsZQwAhc2R/Odso63CZ4L5jimWZ3GSHL1xcNUJWzNE4uLU8bwq+eSN/zM
e0q4LCd0VghzsqcJc9XTaJL0cgm0BkasdcCpqo5Mwhn2dzGJYdXDEAPC9pJivrTgu3negiO9tT60
v0QXif4ZYRaq6Gky+NEgf6ehF7/zlCR14g5GmWfQ8BMOvclepOByixP8MGt4EozYP6JH/ZCwYu0X
Ce3VZ9lJjqp5ymPZ1DHMueO3WnJcVQA2cgLWfNSV2UO/ZN5gP7iKCfJFezok7EYraQqm6D4qm4uF
TGvyPu5oeM9s1YyHJmyF1+GQpr9o87tf1DPrfgyUqPCeqIouRSCJR2Ofmu7J4q9+5vUqxzR8mJri
mHVENeZKBrDqMMma3DrWMHHDn1GmRUmHRruwBahu6WeV6F+xUewk2wudTOZb7XgtfRllCtfnat0T
wXrQ+VNmE4s5Fl0iWHd6eHk6CtoIaywRrFl/MYU/NzI5BLmMlJaelWb4s8H2VPWBr8iVwZlXAcsq
uH/cTrBJD+kwcvaAmXHx3VZvx119uUFDoXgXaChQD0S8/R7Z9NmGl4Z1JXKLx0fhGeAy1HociqoD
jcYxAD1CdbTVqA+neMzfLunkboYsF7uZPD+xUYBICN7Wm+ZuQFY2cUYJ70kAdyHKS2IjYGo3VyDo
57868mF3Luz/8G8Du0biLJAD/ij+pqibRV0OYAWh8NbP2DmXWsC5ciGYmpH08YDKnNreSt3DCfJa
zGAMJS7A3PHFrAuXQakwnMz6x/aOEEFygMBkIWHv5fPgqZ7AkhWQzgO0+ud2+zbxctv7XEj2maHb
qr6dgIPbE3fXKdJM2kmqXsTzFjgvmBQ9wseRlAGVAJXCikEJczR39cfA/W9oEgohCBffmq+sExkn
9J5JQNX30wMj/hMHcVpyzzZiqW7YIOXMddLwp3AsAz3TMyFaz3K7zRjab6PB67jHPFFDopYRIK55
iGAX5g6+9VHoHwE+5IFeAGkGZTuRThOGO1y7EVoXs/EgTXclg4+Uiqk0qsXWLRM49lSF5lTpBkcl
mwzZgju3XjqTOnzAjE+isORwgw2fO/n0T7ihNOmM3+pm/jby2X58bXMlkGkBALXikYqauqu4ffWa
xJLORByvFBD6Og34y1e/BOxHyEwQ9UdvYYbN5WBndCPKEpl0tAWpanJhUAGpzW6LEbOOn5kdsBIr
lYXuChBoQK5zVJMnoBsGrwy8ktz9KRJOzTEajXXsEOyLkUo24jTDBGVGBl5AqnIHAOqyh02lfNJH
oQr7Ya2RdEiD+wQNX5lozit0fnMHhk6aPHDJrxU/8oqG6zXIzk6RuCVnMGdVWRAqd1iPSAXvgFjb
PFhm5gYJLUGo5SwKOBLJ5i6gtxaQQ/MDcP7nHsfZTL1APZ01lTZxElDQpLwpJ8++MJlchj8SULdo
a7II3PL8khrusof7SHQy2W56ingbTntNywUjOM1YHqKpTfMnjS5BA+23yodJbzrikIYAAqpBsobY
y4mVp1SnwYXYXXQswuYwgJ0jkhnU7BKqtEEuhVNM2WNQs06bJBBjZNyDWN+kKsry7eVFhw95Yda9
7r+hhbixRytN4RGBnkVCYxYIfEFLqwEdyw1X4bTAG8XFeTqgXd0AVhc+i+CLI6n/wMT/jB7ISyqX
kUvXRrhWeGJAAFF2Y1sf/zj3G1YjB24UPa2M8HNCCeXIEZh06Su6VTpPQigckPSXCSxUhiDpKiPg
xx8S9PBuFnAog8v4psCABAz162fjcoUXTR+TWNdhjI8zDtx7XVT1sgLW0IEyNessDEc98679untW
hTEPeIh7qTNCBIwGh9PP3MYozPfGl4NbAxysXOEkSPajaJfAQx2f03A52AlQt2oupeNz45x3a+HN
vKhQIIQkQ+qP8H9HjX/Qyp0zyWkDKvfnYmyangIkjI1sGZzyoluRottj5LmUVj/Iq6bVRruUAhko
VQTR9hnMsvYeKIzPF6KLAikLOrBq7/NwfC7CGW6i21NnH3ygaHj/YI4uvh13tzgfvtCts8Lggu4O
4g33RZm/V6LQAGtVRXbTTMpoWsYqlYZ8GPR2kLcGueyC+U0DL3bYFrss7PHdCyCJiDkrF0kBnAiG
C/L7cwbbWq5rQVhaMez2KLG8KoCJuOKERNKFBI0LUdddGldw07wgHb2/qvQ/t9aAJzPfJ9GQwVLk
0PSyJnPeKYHeZ6pIRSPRxMDOI03jItdCofeTPjKJOQ3PrmuAHmBo+vrBNgio1q6HdXS3z6iAIsOO
F1XX/CMJVsy8QHuYxpn/bD08NLia99bThCHNkGn5rJa8CQHu+VFo4AXroRGFEZtcK/izjWoQIqM7
ZCB1eowm37RlQmYP+vysacnKoCKRyC8dqttKD+ynSEBpr578JZpuszwdXIba9brBrnf0DdINE3bN
6hkiKXuFGyAR6iuiE1PDpO8MRc2+asGvPS00UKypFI54cTjls0suA5G3xQSwwYpixGi2vZe4AF4E
+S8j6lXTVDAoRHlUUsOD3OmoojSY1wCYe5/pf9gvSDAvSh7trYwWep/O0FBSQImy4Bo/E4DuD0R+
mWieWxwnW4unAnIMFDP0g91fxqQbRjm16pfrphaBWREQM9KQXnYzu05zCcfiPyW7zYBrOkHI4huN
NHfFQ68O8/ZLN2lRx1d0ukb7NUxkwei/qMXWPiY2iVc0Z3a6r7AbH4wr/ACmHWlgwbSroUT47IQl
feA4wZvBF5RIFfKIzym5zkKUcThH14BS93b7S9RnVsilJjuD+r8aPYWSeeMWuNwuzoswE1gsITEw
vOXpKFGcdeJJTzunvMAvNsfRrCG1UydjQP2AnURG2n9dNmoclkC7nk4itkR1SMdhcmmHWEu1wdBH
LVUMn1M6t6dgQ0Bm8osHqYe5VY8+MiYI5dZ3P4VWLLslZ9+ocHv+vMBfwGl6/ZszgXiMdYXuWNX4
JoLacvNvcx0ZOEJhCZpiLp4H27ExYQnUCTujmcInoH4OQ8lvKyat6+eivMXKVgE1MJ/yGnzzX/tB
Vr5jqvcHIPUlB2az19j8QtGN3n40MbF+CmcB+LVMckGEJPT1eXQOgd3dmFDBDjYXw7B48bGY6Zrz
AkemNKcHHFCLDPvLcAFuvrb0eEA0/wlWRxkCa7ogwPvZz5Ek7kRik2WoKCWY90/VktjPj8nG90er
nmcgIpPIAhCgKrFWW6/jJsH5r3osRYVreINjKDJ6zlddBTfp41TLuNJ8VkkrZJIBxY6jNX9SN68n
3eIZ334B2bbg/9oHSAEKdvzkq7dIcn9e0CO1gr8TyPVMHCGLDWxeF+o4zvhNmIAF8bg5y4qRXupl
dJWfzWvI6tJFdLJycQOjL6wV3D9zWC0uAGtBVP3AuauPqs8u+tNEkGn3VYyMovcWSNI6+3NGiWhm
wIoAshAUAIDOTpL741GV/dYgZZboRxvY34xIBiuFVm70moxGB+t7ldaevysHmB8KibzrsVhKlLJA
5FAJ1EUWdpnluw1kBSJ4qgTggcDE/wmYDM8OXcv3inORMhSoijsQfrYuQyvf8siBN64gmLASQ62u
xazKHLpYDagDtlmwtayIdavKTLl5Glmpae6flKshpbeAgSrpjW8J1d9ro8efgbGeSPmgtnBzclkp
Hp/McujcAJfKL3DnqhEwzXxQoLv7vf8nLTIrJYvjzYF2mhu3KnKDZpWv2h9wGH16n4+o4g84Xl0I
GZ6Xuy0LVWvHldbz9UZtjDXMsDtDvaKcHE+Uf66+/UEMXLNcIaKD1uJlqxQ2JwggPnPtlxwagnbk
XtWt0dQ7NI1sI5DxpHClkFjsSCm2YLMY5Y9iBl4KVLTinKmhc7ZhFwzTUOf/3FwaslEJYfEs5te4
bzZ/UpWW5trf1jiOiRK3w/V5XUJ9tF+gioyYx7uDUptBoo8TSSjwvv4oVm+Gvl6HDfJ7bdjhKDK/
ag1VjCgvIh8xZ7fDSr5m86P80vretE64yVLlwCRAyGwBNY82Y4OUx6icXcQfI0U6BslnwW6OUaTB
qF4GKg6SU6RG6TWycmjK2pseWlz4UpVn6j5ncyKIwIiAJAH0YjEPLNf8Pj5R64NiMYPjJGbxfQIM
EImPnW+KyxjHCuutu3WnOHV4sUwrPez2BnbzUh8jTXjc1CBWckfzK63KZE/OESHhVEEarmq9ldQi
erNW9CCqn8TgF/wzhVGTXpYsRDcofCxUIBzJ4ms3/5zuh9iDjJ/pqdQG97+8/ZIahuNhfR9E6aFn
QtlP9hPQPlY2qOf5AY69j9fsR6oLKK9gHMlNuYRCFWA/TmdzZKHXRHXI0eRKLt+WwDRluXTQu/d8
nuNGpvbdZ1yV9PhNbZ+5ItuDzwRQAcxxYsJCD1lEWPA4/4seruhtHP0kmAbKiROpTcKpQ5vgL1Sy
kKRMf48OvkO5dw/NTqFmFo72S0cAiGT/UQyiNoi+dZpWAstTSSiXZn6okJaIwayJwVad2iYtqZRA
UTd+OnKY444RPoiOyJ0cwQ1ZveoDgnaZm74tRRWffcP3fn/hIyWWWlcUVYMvwBIHfpoOmDJ7K5HE
UbzBJRWtzKtFRJQLVI3d0HABGpZGW+Y/nFgI+6x/gwOixoHSDn401/WohnZp4MXhrkqLqsRW3gHu
e6RSsME8FW3A/5sPU3xHVE1WUgcbK1a4poHrR0r5j/XZt5YG+0ElF6nSXJaKqXQxirmXStH8Mkqe
Gw9XwdMtt6fxKmNNorDadyiRkVxZy3h7netHFbK4VS/492Fq1kthzvPniw5xVjE4V+5L2TgA+6ji
1k0AD3C5GRQkGuce+4FMLhka2BW7srFgxP5nVnfhWb0B2vQeNzwt/FRCbM9PB/bl6pRVm3aZAILS
6DYXTO19oAShHh7RQGDXiRU/BzlRSXGQMFdo51W1lAq6YK3ISOfnmVYVmAMvg5jLjleQSvDEqfR+
vuPJpp0BchYSnkxCLy0baC/Pnh/7+2YjWQFcBulLwoTWSUmXpM19cWcqdcpzi6nVyuavqSrOqWy8
rIcEgQa4o8sllAOpJpzpvk9C1tkgwzrk0GttBjQ+5qpkB2xZ0KmQCHPO9pwG55th+fRceMxH2uMA
yk9iHT2w8MDLJLH3fQ4jd02swpv/fe9QqDxRH5cdysWuAdwwbovtJYHdeSKYnWaAckwINHOG46V7
+B8iPhH1dqjFL/ncRL/4n1JqBSEhmxhaBJxSGcmKbZ8vDY+qo9DRY4s+TjQRVcWlcSHVIZNJx0XZ
Tki0duXUI/IHtW2kSw9DjdI5BwmNrnWrkNtF0R0yM7+j/8iUm6FOs8ffyZVU0Dh7XVnVmwtA+ACx
zvetFFefw5KiOwk98GQ2JnmjoWmmSGig9gPFCmhleCQdi/VzltmIdZjOsR5y/RL8c4WxS5smF+Fr
WR2f6SqkeU4pJ9vEVG4ctR8eOqvRMiAPGfzDOpO6jRuX7QwlGwaCWZLv/cUun9WrUqVQSN3vp0ls
j+H+yDak8EvzyBbREMs3c8VNowL3yX1onKU1IjwQdHTyv5IXTHwLhvyaM8/IV2/wcN8mATJquAzx
LPcEHq6ToM7MsEZjgZatZGiYgERIC9B36UDPdXcSbfEGj1B8v6co+AP7Y5uJZ1zxCE4nQ2HEZ9iG
Mwoc+eHDoKqCQZZ0xngJt6D/GMAd9QVwVsUdecaNy8K+9hruLkKspU45EH2co407iPWVZevAxGwk
lB+ZEHvyL4rWT6VBJiHYGR35+lGiHwvrdPisMs4OvvqmPWLr/+3mopopgoqT9JM2mrfmHrTKwFfT
xKJ0W5kpAeQLvjkaA+aOcvtIAykxqPMhF7PHUSpzUd+/0n0oEMzRgr063zQTwV9fsmtpnmyOvV2h
Czg7Muqfdvg9lZt2Q+U6gvCjbiFUVytO0+B5EN1LEfFWMCH+R/UB6UPoWMLBXD52HAOhA0JDbGdx
JsphLoJMQervzpqd3amL4mx81FcChtzWX+sO+GqvXU73kRwuS1Cvfyu78H7t5DU7kdvIzqlu82Qq
owUNJ/bXRSZmNkdwcrb+UjN06RiBN9BebiZw4yAcDPJlUTQhXK00/vLPugTK89A557BO8Zm+yGFB
bbApJVNUF4xBaDnn69gJRNmpT6PWGaO+7019ujnXXUCJsQmuJS4/yo11snkK8AxIOjj0/gBJU2cJ
s0xxVlIom0ZWCOYSXp0cR/Hp1Mzv/fQT3Blr9Aszqgv/matnt4osNe9iTotRlOFnIF805TbjeIjF
S0bjxyhkcgASrje7n3TZ69QWhZzsNeewtH7Q522jmABQnOlObt5Z/SdXrtWymd6Q+k3WlafjCnuS
GEzM/Hn/1Jv5C31b6E7UwAMYjqtADzAFZqCAeAz8tUS1j46HxnN+dq6fubYafT9VMC+OJ/NxcWHl
Dt00XTc5vVH7MjLNLOmAgJMoguqcoN+2RFqfdlXqRiZxAQyRoKNSldyeRFXwvwLQK0ZHwBa5A7yB
x1ogMVCbMCciiBSRGlBA01Mec4jj7z9erJh5f/BkxGq+lm7gPMKUyWaz+LhTeYTYRpUT6pRUWS9U
ZvA6HOvFuBg8ICgmeaU1G6C1vI1gnBGsT+nCSqW67MH90igOB0Urs1bsZJq0Jsj37hbdcRvBkNyX
PTM8IEC2du+ZloZMSrY2lBMAvjKKTNlg41G9O2/Ce+iKZjVFX78Pl3YBIaH8gXPvwwzsJJxijjjg
LLqlqg2yIOOCZ+IERtpPeVCVdyYR8A6HVNhX6+tGTLljrLP3ESbkBnDslz5UiUTNEnYYuSY5LhVB
n+oUE5vmsWb7zSsv31acIQAX4okdz7dQgsVG2JVqrrOiRla6P/IKDS853od13+tzdimn/z2HmVik
8AAAYlXluj7Grx/f5CP9K1G5VPfUzx71rKDa74Zko0VVDggX03LHNxoRdzzLt47xTpkANNt66ROQ
EMmHoe4pRCAJ/xv1IQjeof3qs9fHuTqu7VaN2+xruz6YHq4YFJYeFP0sCa/ooK2S83joa+YUtIhz
4tQgFc2XUiukHlIyspJdnCjp87/YFqAKtwthnx1N2I04fF1xCr06JmJ+wjxKoigzVlE2GadzQzzW
/yPZKzD6GE6cpHQmeGoU90pDGnAbO/sjXL308qJIDuKuOqvDax6MZYLwP76l0t/vMpllOqbyxQFe
ViYD647FfJsur96lAvG9oqN8VE6k8/mN/awgO3RqHjzqK3JwJY3ZPr74YgRa5S14w/QmEnq9zqP8
wOtQL+0K0AyZlKvcSBJHHjbP3uBO990s98S+UU0KgFkQLagmdJcx6RS95B5uF4Ze34+6N6oQjGZ3
t9qE6Es8MR9FCQCCWRgWUa7qL/bFR3yBGgj+ZKfHYx2FZ43I/uWOygyvmecVB16mS3VKAXZqBTLP
e80VdIo9+IUXbxm3w580yWmMaJPlw7CXGl6ajnNpGYNWZsqTcWhrB29ex4CChLkVOI52+K14+W3T
RceIe4J/Ck7Onm65b0PHe8xioLOez5y945UzKpZ93PLLpsBPfZESaMV/fpB/7c1aA1u+vRybZE0G
1tKTjiosCQ5omQ4eiykwhBfuPyj7qalNjOQ5JDIqxzmL1WFelaW1DJzhI1+MN63+CZoDxEP37zJ8
pT6smeezDb+nFF3j0Tcr+Iu44cQsnIHZ3jf7iDbhpWC0TF03uqn0LFqKlycZBoEBKlwnS0NPiXiB
WuSkd2J6QA6Kvxwrx8HPwgkKURj/PYvpC2cJtxo3FmZEl1xOx3qULLM0c5xdLcM7adXFOiL/5cFe
RDJpydCju7PQf+SWi0NjW8F3amFwIGJmYKr2/q7coi4WxTqutbI+aEjdCLsYtAgJPau3QE60LbBD
fjOneAacNOr+P8XYN/YRTGbxArVt9uvDAgPFfVbFUNqOllLRgDZf4rWSovLpK+wr1pbRuRL4FkRG
impSdSQT0V3D4NfyuLOGASpE//sF3AtZrRwk9qMojjgXv8gBIT+ipf9Tuu9rEgplZBfjOMpSau8r
tRl8IC9E5fPpszeotsj5mRwYU2PKJZRolGySu/dpd/mZRUcErj6xMfRxvqiLW34/UfUfGuQhpf4L
yuPogaYLuZU+5w3Ve/IDJtjXazkghmA5jaKZOqrvst/K0dvlKK1RqefV/l/sxyT4NhwJRQCt7oT7
fkLvwAF2+0rkfnFFnxA5rqFKWdwRPwwwpaJo5WtpUPlU8lX39QLt5QRzrW5dRFvWv0WOT8cMlT/x
EfZRJHyvHqJgBY9s5mbodEu+Q/AVaS7R3RSMfxup/GYgMzMwdgF1tqp99tLfZkNYZTsaz0+zLJkt
3angB2ky4l9SsTF4csHsZ/7uXrG2rOKKirrhrAmC+hMJtG034xNFEI4+DDmN5LVeZd4DI1imaBXb
Jphl8jbZP+kFuB9UbWvF6nEgnVq3HEc9o5d8Q+Tj9HOtXfYbtQR+oOqo61GFgHL741YB6BAxDs0o
vovulNgAhjbBV3CwzDrxA0VfrXwFMgZ7jucAxKsKxfF7flzGSEi+t8kT+FNfpxjZEpO5RX/zRw2F
pm3yodFnmc8N30JTLrl8uQMvHEhV1gmr+SKgvieDtgJAdLI98gbUqx8feR61mS+R81G/ovFtDXRl
Jqx6FupZfoaxjQoUf/k6PAhF2oZWIU5MpPw2WMvXjPB7GARb4kOXqWfF0SNunmW4qsiSswfC30ur
J7+3j8pP8fk83gqIqEBGw9gC/o7tVZx2nRQCfrDuY/hKQwHZeWj0S+hJdRfm3OU9wDWPxbagooEj
6TXmcbQ/AlVPNSCoELQFsydD5En40GgTbIRe+Xf8Snu2f9/tHSVQhFmaEDSs/+gHrAAWdGOb1aT9
uYzpcDw0Jy7iX1awlhbsFAu0CeHH1gJcyq+T4MgGMTGDXYunTIP29bi0mj02M3qLtfB200327qZT
hpSh68yK8n3QDTQGhH1k/ymdjvRcfAn1VwymC2/sL3GIRDkWI34qucK0XTgaYkDLJdPJOvPqoey8
S0wFeR9qywo7CT2ep8X5LsvZBWd3YH5HzruC3ZNRVWIlI5lJcWVm2P6LBxnrgXxdX5Or0emFce4R
G12x1bibBpzYeo9SBu80kJ5sRhBhOW96UmSn192mRUfogb9fjEj4gftSme8fZItU7ZSKGGl3n1OX
Sk7lai67iPlyfN/y8uEU0my3ZgWmb0S6qV38+U9TsC2dxw1pUsOc6RllgISnNgqwUBuWabtKWNwu
PUkPuFx0tyBFbcK18O3JLny8b44NKy+Q8mgiS4jRi07hJgq+V3wBMp2NYJ1ZSWVdfaeHksIZ7Jlg
DjRbxKtwe/F+UwVCgTAhVPHNpmLhkCOtexwypItdWaLVeJQcjDG/W/5dc+O84nDGk/su7yzen2uz
uDT1Q5u0iaBD979vR/QtylyEJ9+EYiaxjX4gx7HuN7KpvBbZ37sUQEZkllOl46wylcP8TROuP8z8
t2BntMF53TZzZMLLtkL06REr8okhvBOvNx381kp/Q+sMgQoB8N2iGI94s8mmfhpEw+VHszQ/rdXq
E//Q4wyNTxm+S02Auy5LXwefZb4547xiQ/+QvfUooz7rwQQNfn/OoMpvSWO+eglHVOhr5Ix7Jofx
Ixmt4ekj5f2I8RY/jsS6FXb5Ve7gc3iEOonmbvbpuVbUO8TqKKanFcxXluYd11qANxiGA+LWmHhK
yCsrWH/dOgF26/qrMDED7wgKy2tqOqezbVuj6ua2P9aZkukB0pqcwo8WU1Xq0qKOU97Hh/4Q5Wz2
hrZvDLVzZ3svldBFN9PbUQumIhCmxfg0tOHYcrghq+DU99ZcJIy1E1Yyfxm6hUp1r1ZC4SlbQmbT
gdOFC/3nrOyvV9khoyl9g6/+pmi4Rt4GEZoDUJJDtfdiHh1CwVTDjiK+5wdGy+Fo887Y+1qHmywO
E7xxp8u0IspirPJNxzKf7SPfKmaOYOiowoG6a9Fo38+LEaIScLuj4ZkUveFh7rWNtyWy2cCUG7bQ
IHh2/eA0+riGnupy37ah1l4Zu4emXqe0Vec6Ax6daT4uGjTH6ncQIkCYY9ws41kpPGHhYdZZgbEw
PehTJ8Q9/MBw+8DDo9gWCTAGpuiWekJ4sM+ywI02aMrtKZS/uy/ckLub1b+8ivoxI+Y0FOftg8fZ
iSzixywFsuztVr3dAwKDMERAXUVu6rOaIy9c1X8Peb0vebwOMoY+5di+BQTCcAQTyLdQYGLO1gjn
B0VSw9bEznOax9/9Hc6Elixgi/VDXRKfu8ppMYDNubYLXLV5saTRlR/naNFt3SH8D5tlt4DzYbaF
6VrdYUU6t6ePqii/ZOQSkoXqP27HBAUPIR8+mn1CMTxe0fCKAVI7R1syExMeDy4wilZLbXs9MdCr
dxLnYDAA4E7wwEAmQ0Ds3QOeEVrOIulTbw3+Aj2jqteXvxsX+6KKJHFp/y7k6+CNYg+g8f53XglR
T85W9HG/63dIiWbZ7EJVHRJjO3cqhXGV6VaBs0iYxc0of4HAauBhtkuvZwYc3LzIFVDhDIbgx5ih
Tkz6H1flAiad4wr0/lgzWvFG+i36poGXd/yUfP6crJODPdirYCVIQR431/mL0qNr9I4/bP4qaias
abcwk82OKCTajWJLWIYEMxlV2422mwWlGRrml2f3VcBMZI0tSKGWFH5UncNTAIWgw2N92qyl+0oM
cOTJQ9pLuUl4qT63I3wAMqCT35/XzfPnVOR8kLICxFIPNt2hrhtfqOvFFPfuzz3JySQhR1QJu865
6C4yfDHzMbgRGTa1iH8iqefePHN1Du3cwsD3dBgqLw33+WSr3rAfhvtonhBtFJVvM8acVoJsRTx3
k5ceqRChAc9sQ6HiZJZqDXZZrYeQWGecBZKhu82YKtmqgA3HafzGWc9zhmIpq/2V2lIVm69kco4N
QSSBS8qgJiqqA2d8pVzXZp6/jd3jf6/euR0kyVmlRdMmNhW9n7eYk4IS8bkNkc2DG8VniU9AzwUy
XF3CXnrmiBnQJPwgIlOCcV0yEjgzwfVZBQmO59dTTAAr5ch4fG16qUu4+bTfAkop9L2oxrVipBPv
D4FlCXmcmxrWriQ6EWPnMhLHF694DCOPMJLvuBtPdc72EoBuGtGbnV6etJG323xuCpzkhLPVWB18
ysDiaGqxOV2vQWSHwsFfpAPJLmrxtZ+dkdgsWBqycJk9tXxvH5BQU5hy95fMelhAlng+7vimUcGM
vm4GTN8h4atzS32sKuiwBlREEkppku0afZqD4ajR2ElqHkfu2A70oiyyyqcn/PeE8i3CEKOrRVvD
MzamzI3s/gzods89T5KKNoEJV158Q9/aqTT4YVvoqegX4gJlLOlZQ9zlqDxL6J62U0AKcPoidjEI
EwVEZfZik/NKN2Hx4qQwNUumbx91wUq+YWAxeM5WfT6o7Ic/Ti9WAjmmXyYbEbPmXE9+2NODdb0r
gVHJBQ4IwFjbfM0IEdnarUpTQ9dgFk8KEByANJfuUBiqFCkLXjRKe0wZS1hEYOZVJyLzRvKvtS0u
TiqrkfZ+GOJ6Kdz93p+zj9nCzA5IzvuXkmeIxOqfICvbcv6IFyBQmVqePDCaIMyHbmlBu4wRxerv
99DBc7TB7nWByMshq7uYgr3QrlM0zZfpxIDoClot6OCJlJ0Ozu4W+gB6mudOxAsQSK6GE23uTs8G
ociXyyCEaPCKWlaTkmKdRvg6lA5fReun8Oupr63XckvZzE0EPzqJ/l65E9Fgj4sxlF7QqdKq1BoW
xx70Yxht8bb9aoSOr0ViTjfDZQgY0hhifIKZex5mq7bvuh2+0CbGsO1jhdPGE4juqWjYaoPPQsaD
lQKobrl02R65AAegT6ETXkP+pi/1yE4K5amm52bmONbKfTxbI34jAA73azdSazpjY/GO1mJwKQoS
GLjYpAIxIGWjn9Z6G2PzjP78BTrwXn0xviU6VKc+kqjpWZjwh4nhNb/1kKmQ62Jchi5xXWhMnY3Z
SCNuVmuFDE7r05sgsFlx7vCoMALR67SC0iQGkw44QjxKH9pE4Ear6gESzUskK6FM+v6UtUT2rWvd
qmm1fjpPTJEKw4bqYXCKcETQN0aanTDV6PZHLJR9IND2Cn9CQDLU4e1Fl1v9NC28OkwYNuiibn+h
tGXCwZpc8+rHqkUR10L5Ozm9gCRVzZGwelOHpZ/GdvUMYWamJHeJShb1tXeKenfgrymMnh6xSPb3
tumSts/MghSfaAizqPwfFjZWDd0kFPl504usdof9aFeA0HU+0zRF4EKwB40dQafP1Xh7Kxjnri57
O8eL02njBhihz2vw3+w7ROE3QiITTvDcEhj65eM4IOuvk47Q0Qrl5uX4hiRNyMtFRNrSmrubquT0
3ubFjHpPPU0FutlxA4WDGsaEW1yHYNd2dYMXYMXxhKKrkzn64NM+uDJTM6CZm9Eie6grUfRt7S3P
ayGC4iwkihkYIAmtZYkYkaHQYpFEAEDHtkptJJuYiFaTUqB+VL9Nv8QwRuoxcO0T1Zs9/ZKUGzrn
wq+TbwWCTQPbfCOxApuoqzpkKSXYyls3gBAhjkIP4Fv4Gp0TQ6V5Zt/EeGqnWnX6HlQ32byYW1VS
fj6FrDiqXW6pLLlfYQUiS9OjgEflrlimYSqm3tnkm6ph+rC8ORzKq2MHwqvHQQjcGYMfLJNIkedN
pp5tEEJf5HAfUfPF3js7alHodgxmYY8ISrv2X4pIOfrGupfdrMXEo2/ct4MRrCOTbb4iXXWd/eHe
RlUC+zi1EKEvkSUV2brLkSnbiPEqTCtwqDGHA7nEt3v7TDB/f7XeIykUWlcsp3sah8OMeNqWpt2Z
d+AHktFSQ6xzOKhOoPAO0SQ0s1zRWO30Q5Yh4F5AuQatTSp1zUCcyQUlF1fvlYA09BJwpdQrgaMe
agnRvhPyB/aeT7MPrP5xdJcgH9fzuBvVn+c+R/1Qal7ONCk6Zkop6O7bz9ZlxIULtvaUMbCfEtXQ
PXIkBcXVQLx4Gn0wlvOb+fSSPYInut18mYeztIjPAhAF0lMyE/ijMa8qi11TWUz5YNWhJUP5pSrQ
IkQmZIeQNOWtYtejKue+2m8mFnVAHptBcwH4YD9VeLtDQohuqeB1kSjLiwtXX82HsnxJATrEKhHF
CjrYUivdzxX11p6KqDBbd/D40pev/5YO3+hsfU7/MLLaqNJdAbwHhocm8cgODWn8BODlyuzwn3US
O2yfYAK0bVsL05oT4OcCHSJ6GjWgVJbGxcLfpDk5Pcmwc1+cUw8wzpKAaq2xipKjzPya5ejeR82z
6B0cNwVNrvrNUPfjw3BvRua3sdyYKjOiqkTTv4+MByvOZGUfRnWpzzxPbR3KwNCWdVg80SB9E3G9
fq8rJfr2P+o/MenebONEEwuUN4XoSWSaS5Qljzn7sF8NS29uWThbvVfsKbRqdqQwxJ3hHWm+QzsX
QwXE2wok5LQhL6dX8/4sKntAU3OVPN7fTGoSA6GX/FnLnhIK1G5rQxWuQ8hVHnARWLZUIRT6XREw
IZfKCeYfQM4TEM1ReYZzh29Db3Vmj5FXR/kFKB4qszFIR6ybmtfsB2TwH7aybaWsO84RmJ9lfWHD
ov2gLcz6Y71jVJocdkRouFa2dTr7xGs0dXQHhM6hPK3eHDRcafXlYFxz9Hio7CuvNVwHKiTJCFBE
0ZIDQNmH/741dRsNeR+KSRNZkSEB/C1tHleVm9iKgQrRBbVNVTBqfr1fwf5aH5R0G7pOWKDyUKwR
MVs6p3znPkzVRzfWg2uvqKMHryqWBiVjQcbZIOegvKymi+asOr28jUdZ161Zq0raLXJQwXxCSE7s
p7eo+AMF5VMZGHefcjeZFNoF5CyVtgyjtfBN/EZekDEb4YPH7PSqBHLWJxMSUBrqvjsXJK198Dxx
TbjiVK2EQDvCxpzOw4ZH7NhAalGUNn6w4PhfoalHqfdRsZqJ7VI0OMNMCr77RKqPrRIn3c2uHYi3
YTjtUxm3jIdGbBRfk4eJASW4xFUDZfJffDrO2YZSaVbuCDpG/3+JSYmQv0FVx4mNLvoF3n+8JsJB
dqcs078pSb1Ps2WrBVXIVjMOJ27aavjjzBL3Vn6gFyoeoyt2Ud1ACiJz4rvekaareHZbRKZl4i97
d3SKjkzwFtQNtBclr6GP4ROVsGhVzyi4qcjmQD0CLFwILWY8brkM4p0KRM5JnN2qQhFXmOgGGQBR
14CVIJRvw1dmMhRigDfByIDNxhFor8hHe0gHjFM1TjlcQaIMdGiIi5ZY4kivbNZJwDpZW9ZxPqWx
WSTCRXWc8agiYHePLkcBJt+KUkyCK/TfF0sQhFnVXMnoMi16MtOghFOZvkGXW2MaJjycOWhjjiRx
JSwZ3EmORBWJiktlpdcLaWXKYl5HFEpMf3DuD9DHZTEU3578PdGABgkFZXokMbElYeKg2HBli6BG
wWCYWh1c6N4OJzaRoZpuYV4om1hre5sXPZjj0/8XFHAPwkNR0mJ9F1zBB0X5X+uqGufLYivbyddz
15oyC/os4LyR2kWXsQ/NVL/XVU0arp6xj/t5xgFezmfvtieo172q1QSvE+ASgItDekzwpxs6gONp
c62dKdW+v8UjJqeLalwRHny7QeAWnZiDMNW15UXs2+eMeR4YbWcXlptj6Im6zUnhY9N1hKAczyp8
YTxXlVJLEuDT3r6TSkDlIVQIBTXLOiylmdosV1vzYKMUFZ+X5BcifHOjP9zi6ABRl5kceTXA+MRt
Fl9MavyxE6D0jw04q6n8RI3bPpnHrtYNS5jsT7wCY72MkI82Zie/GCXs1QS4j3XaEJgZsZqiXU4L
NKfxhuyThblMDTfYCFqBavg9uS8sbOTUkJMsyKBnPjjeCTBp6QPUILRZZLOEEBMi3naANRG0Z2gW
p6v6u0GPTg64Qxxen72e65s4I6qf+gI6901x7MDREQ6lyjT2MQLiky5Xsh3NWPFan/tw8/4tQGbk
4slL9qqIPG1TfQg5QTzJ7Mst+4ee+JBNyR2Gg8idC61UDAXs8oYkR6UaDMUuoNmWD2S/mm3+QZ52
mBoioxkXoOFepZ0XN55LRZZZB5f/nbB3fj9skfsQZvl0do1RLEKT6tMCYdHii89nWIYbxZfoO5aW
Oky4MLJsQ6ov9UOLd/wwz+j1ZViZqe63UPIpQ99LzXcvt5FrCm02BAJsHrmfETX8ThhWxXWaEzSs
d3l/dgY3BGs96aF9IKSq6OTbshlzTrGff6M4T9kU8JBaZFvu77TNbsT82PtcOGbf9u8Gv92cpCEA
TF5wVgIE6Qgv/XaqvNH3bkNE7uE+UbUoPJNR/uQZR5fQVHpUSooHXmdkExIUQYaE2OAeut4QDVgh
oSTmy2YsLijeI6E1q8KU/jyjAVREpYAvCmOQTVsIMO9EmUwZjDK4kWDceJrofjIiEOL3G/2WRpv5
sG9LIEehsoJ2oaLmef/C77Szpmt1HEAGQJDhW1VS+GQdufagbrXJqwp3VFUX/ENOBGZo1JZO21ag
pbqkfqciGMittXcHxCHYDwjpdOBQUQAiOvCv0tMXrG61TFiX/3mieOJeTHRIQuLS9oJwEHcfMTE+
LCENGjS1ZaSi94Y1SNrdCDozAbQxRTvufxj/ezy7mK9yLRLYkGtS4P0PWV4A6pNOxAW8xaSsBedt
QhBmGZmuTk6aPdJ6ZqwslNWe5/dA+H5Gj0Ahhr+KyVYxAvtTz8/PluhEUOmHqjDXgVtXu9Y1O8JD
CQ78qs7r6RMZ/zrkEKhH4vMViMUI1A9ToWmyslmtcS0BoS91WBqStA+gyK6eSLzx7QEhf5m8NMOE
h3vCFnSmsTecdbR8cVKzGla++7BN7KahiIttaFc/pOoQ6UZmJI/0r8psln+sFxwzb4jpMPeYMeB2
EzDqRvDvk+0KR29XxMWUib8nIKX663xtpAnqWe2fq+/2CSyAFfNHoVILsAuw3njt97E7UwEogber
1ToSrKLMAbnDDXJQY6iqLC6ojAJiV3txxDmOVjRJpklgG0XE9uYlQbwxVX0E7svbl6DOB01wYgWf
rZhPPFDT8CmHQRFddMW4ldLfhfMX3AnOAPAGi3EvFQcBf0GDR6sg5yD1YkQIGlBa9vzEBMz9Ng4B
8bxdYMPmlr5Bc1jpHfyq0NJSblGYnfrrbu4lXiammOFK0FsTo+7dM7MKMsllKU616jXJpw7NEyvC
ZFMQRi/n2C6CI/H398yszJm11ZgYrYgb/3ztdn+I8bK0UiIuneUVKYb2lWFcSS2ZSOzRMBOfQxh6
mjmJB33vB8pPGhLW9t2RLbwLK9LDF/uJ0AWx/unmcIJ6pTgqDtDlA6htXIsE3y6Yv+klT1fNvw7Z
QAXnFmbx9YQHtGzVSF0+jVhbg29TwavGrKh+ak+RQY4S6CI/gZtOuCgumXuQp+HgQwy/JNN+wCMW
8hbcJWI4TE9PjyRnDb+dbEGmB0lIjIDtHO04MaRu462VIKpM6L0DK7uh8AIZHt+XJNkWjTqk9xWE
u8Z1YGZrBFI27G6NOboZcYs3YSwkszM98jBrTbxk4r+zd9rLjbIzdpSojq5q5hQBbee0pp6JjslB
wUHnJr0KlMBoFQcBb/ScIpW15OyL2WuWvbxEKH2QKwrqBk8xymbJPM8KAjxxGUUd/wQkzPfIrRGn
DWDZRkvAHhwV2/5vTLL+TNPRsoU8OJxdoaV5g07DJuwoe1aa4wY3cOlWOB2y3MqcIEGKKn5HZ24T
IUBiMaraNfZtoR9MTEBjq9d0j/rYjzoNh0MH4SjyKnBwfhzp5a+hkN+DEWDPFGGXPrsByQ003Bra
sBGJ96le3+KtWAfVW4KxRJBMwGbZ9RbSAZB7/VOGWSC3QcejV/jdsy6xaVRvikc+aMVRf6D52wgf
g6bx+QtZa46+uTfwgxtZnkrUV7rcIYZBLyj7IwLv1x5zaVfJc8NLc4zA57nx3ZT1tHKV9W3Fjj4Z
nkwhHi6D5sWgHCQtHu0m7QDkW3d3I9gjgrFI8toA6JOHW0BDabBJ30Qfip9pGz8Hl3XAy59ieP1X
3MJ2p+muU/JFCtRPZVQmVydf5sWPNM0k8byI5qdgT2jDGLHmtaS+mUbh18xNtEcGkq5cXQdJeDIn
EvX2Mx1Dpzc8TVDblmPHW+Q1PiG44VCunGHjYjPOvrO4FHKUcu5rNZTNp+VKMB/95vDSPqkpvCOz
JeE7c82lv1YXY+leR6OXNCn1W2IHmvsiZ3K5CdwXU6ivmg48CxfoXn6M1sjHEiA6aYmpUjb74NfM
jz0uzHpI7NIC7vspNjJwNXlGh5fgk9aXAtCM8wHZ/ExUFoHmX+5EnVpPhzMl7BcBYvNsdK4YZ46p
yg3SYei7Lo0Lq6HhFW1tzX7c1Dz9yzex+x3qr+1GOCP8XCizqmfqrdHqO9pbVTT7btm+ICB1um2K
3yJgvCJ5lqO9Xu42sx2WEti8Ag/H0+F3Z/MQSxW0HdM7Veb1GTtu8Z5k4JNR7kMwGjlI7wPNJZua
1GAGEESKUJEeDcPXYZyp7D7lFW58jTaZ0cEF7ipJXqM0WdQ+wbEvAEjkAlyHB5KplBZyD0jouZ/q
D/NHII/EBAJ+qOB5rHnBWymQuwUW/x3XQgjcPlhMGHsXpKBZL+ONd7yf2hsEFsljZN+het+x68uQ
ghgUOvWgAzG973RX3DbMRv0htRM25PMD27jZVDzhpA9uWKB+MYAmlRK/0Ch3ZZfedVNq7VKPLy8T
W2/X+f/pB0QPybcDV8qMqfIlWpLeMGkhsyT40cUsMd1lB7eFGZNI+2BXrO5MtIIY5aPGH+Mb2SrM
MSvxOZC0H9wffINblcz89Ax1Of90Fdr+2x30kE6mQoEq25QVQlo5dMGv8vyFymtFnAanlh43yG79
h8pGc8T1h9Yb0TW4i1QtkH3A0O6sGBzCGG2XBX3s38V4rREuTat4TOa3rzvRqp4/4UlCz5v3SeTj
FoYAzbXaMLmJWioU0TXqxszrBfxJrQJGA4hLF4B1+Spv7GuX7PeDDD0uMom9qt99ELZYDkpFPv2R
iAevJ0bs+hgR51RJsHZ1nmyu4RHNcpY0AYHarD5cTASvTITz1FTNbJ091EUF9J53EzlpHEI+Kg/M
T7+uNGTFicrVaGNJN7lL9VGr8tGADpvS+HrU4bO1JCBmapE/nq40k9z8FdNuI53NYgQiuWmuAmsF
N4+Kl+vl0jefpeODI9J+bXVDgK+IjvlOTXYcv3/AmdKiwJqORS4i1uukofEd15oggOuczM4cDTdz
liB3c5Kv1F41+ij8yi1bgANv+fKQcpuk/tb2V9n7nnb3Kccid1l33zUFnzH2KkcHz2Wd+z92GX3P
Sq2JvWNZMrLSaxRpAcmASFZOfGfD9Z6L85Bs7NgjJ3nh74DaA/JEPnhGpf3Rv49lvwRuSLyu21Qc
HuNxSUVr27aoczGmk2Gr88lXDf2Wj3RybSQ3kipKmBzspwzlrRsPRGerWo0ckq8OTCbRGlDVWVBO
rJGQrdzgp6R6JxnHB65T6CkCqQbAbSN3tnEVBKlFEkwCBfEkc3AHo8c9ST9QXyyCVu1jrdvU85mm
WgO6PMRLC5dZp3tu+uXX1pOZQOBRm3r/c8m6nKs+e517z89A3nDkckc1UHM1hjA0bOokO4rHx1po
UTjvXZNYwAi17qD8sXYXR6Aoj5aiT9Wm3GAvBEmE0W+bMI40qQoFoxTh7T5AqYMNZKhia7MiE6h0
CSUEbHnowGn2UfaCrmoQhicFVt6qTFmybh8SFuj2bxuDQ6vqj1x3XPrSsfnLsJlTUjAENJM64MfM
oatv+6mMsfnlHFI4LM2v1V6BopjfaXcZp1M6U8Q+UVCkhoZes4yiXy7FwTWITLlGh/WWhca2v5MP
QNbgsDg1bajBWzD1gMf2AH3aCnG9ZB+2rWzHtEZxBDcb2JX7tvX0dILcGgNjJd/G1Isj0vnXL0WJ
fO90k/9ZC7lTVz0GgrmjbEET5tseBAex+ZtdNeZDN9diV87d5SlAlDfdgz3ORkIPj+F/4dbzX1a4
BUxfN91fel5R8yjg9C/LecuUDbtw/WMj4EJtVu5MeWPpqOxMNQiS4DV00j9akBYvWS44Npgqv69D
CmwL6iXJu4UnDYa8JRoCjdVd+1jXEwCeen3TZdZ5gM7+akYEP+wIknBxwnZgoVQ7gX1FGOX9JZTV
Kc7yugm+TL4vzg0xRH9nBJ6MU4DrIuu8NcVf8j9EZA7Db0jwJwDm6cE2HupWgEOGai1lqj9wKNSn
X6mrk2VM3yujL0H4XqoXRa5RoNzfkgXbroVR+/tUcg5CuHeao/bGcyz9/d9hhPkpufjwO+11gMBr
bQSEIYjH94HYaCbovaBHnGdZJozrZ2qtC0S6Qd5FkUrhw+nDelQpcvWHjlfH7jHTFqkTAtQB89kP
Am/484eoRXzZ9f2InUMLSjcrQJu32VvF9cNHFTuLaq/4XJKVjeniEoAu5rVvJHXEdgDpfpGwZSDf
s+armd/hTgk0GvONrglVkbBrJm6WaD5X6W1cXSBT3M3Ckvv1Hbta5HAO4OLf+HW0RTtXZ5kZ4EwW
xr4pavRIO0bMdOa8mN0jYSbP3PewK1YyBVTa9rDz0jXFmGtSFkf/xFFrGRRhfMKDnRriFmbgCMFv
ZhQUqLzDe8DVZMchGamu3OHeL7hLNyKiR437lIPPt3FMKMswb7nboDL3SbThJnX71eAuv+b3yUG1
eK2Xk5IAeMgzawbROn1uF3yUbT8qBDqgP93AbjsvlvpatP0mb3u0PzWxLajo9J3hDwVqMr6pE+qh
WNmxEaDzEwQXAz71yC7EXujRPcbRsChnJf7xU+X0rE6FQnn2KKOKTVMHi40XlMURgN6MqeCFUrE1
xKXAY9Issdz9FilUPJj3f+HNiIwrJWM7hW8ZTsFx7feR78yOBuVZ8Km8b4/cXulIkcVwPVOHo3+X
bwwu4Lx7f/uRO9k6OoMIULSkdmKL1FEzsnGQwSzt2FV1t0/a4WCoBr2jOqaF7/jR+oc3MH6tcIl7
l8asK9UVSvXgcPAybiPSSmuueGlJLPMJJYbCzd8kwD0g5ic5uNVocFC11JPwtfyPL9nAsSqSci20
Uum2UMx5HuTv9f9ZasoL9bKn2sBYM/YfZpSCYBj5QKYzXF6sD6SC6+00y+dvme8xUuC3pY3bBaan
1YOxGhSiLH3tJO9KHO7uisLJMx4v7MaGkt2XL4LZrvfr/imkPemjHgVcUnGbI8u0pV4A2jYPKpRV
IWdWKMM9xVoQ36T84NmUESYpxcpU97KfXMfn57tMT+HC1ZXF5iVQoTC04ZRvTeotaaEmZOnLxnP3
3mlZHoGaWfk5+j7y+cxlzVGl9aMAH8qVL8YVUVM9BBTmnOi7vhRy7DlWryXqnqMQSJdlZdPIfmrV
pBdKHbi5pfU5jHjmB6haf9WGJxgzS6h49yut5iHZ4WTdh+XFXOvrp5DjKsZ2Mi9KrTRy30dYdR7Y
r3PxQHscUFFTRKCBVDp29+CD/fBlkpOFdcttja0SmTQ72oX42q0WFhy323tkV8h3P/KFf/NTMLPn
nVvl4e4VP83Bk+X861swJDIc1TNw10STOAuyLQN6VZ4rscJwiV86sQlXUyz15Cw9eevn7eqX6NuR
83mJ7+uP+59RTd1ihuJqDRzKBO/F079fvSEAitc4yCXFRhAa8H9hRVFl2wYbFjU/8KkC4NpHDsRW
vVGE6XFC7RHjFA/Q45k4MARqAKknZm0Q+6pXHXBm5JjszL/wPN9R6RGAiMeaACqa4uYVPpaBtIfp
T5XOCEV74MR6YrMQllfv4Ndk+K0QJlmOhO+F3K3HyZWn2lKd4HSnMoptKWVAJtN47+K9za9NBXAR
Z9DHQs5q4ERA4NdIFXbvFGAKVrM5ac+fQFwZSoV7C22K60hD7+L3BossXnfiKPKIeSi4yo5OddK7
N1l3mse1dkeSp02fdcrAlZi89AXpRhs6jq/01i5NUhkwiNjuI4SqqKR8iqKeb3ukDS/mWK2hsJJj
rG654xc3i56s63xDlSuZ97PH72+liPEJfNZxMF0BjbF1aAYTLulTPYJ2Pg+g17vxHbkYxWHPe6Ds
tvBbsPnhiWaTGf9mKPd7tBTlGCXzD4NZIoJBC1vgGBoQI58Ir9If+Z/ol4xS5POt2amgwfke2OCk
mG7qfCoIsc4FeYVtOJFUfijfNN4EBDk/l1LEZTchDkoucPvnq4Lxn4+b2pTUe1bE2Uf5djo/DMM/
nMyAJttWVUwgBFk5XEKDZ7DHy3HNqFjHaR/cw5NAi7oZTB//Yth+wGuDSF+L/X/vSeQw8ri/Mume
F/9j8FKTkUDGriuBCm39iA2TWzjxIoahe0q0egc3VNzBfM6AR2/V6P8681a6Z94lucyok2vcHOUq
Rq/JS2I9tpUB5S6EQWFTDRT992K4x57PM7haQPq7B5DfM8C/Y3XsInMgghVmH5NS7jBUmuQQ8LTv
zSiLWw88/Jve8oc8Q0DOR73v/JkCd4jRt2vdouAmvNMsCRE6LXf0u/gHwB8WKMVmHHRvRMl0R65l
0XijBe2ubmCvAtDlAi8jRafvlpV4E0ALHg3+EACKpmLjopg03NjLT/0CKsZMHojMQ0cZUuWaqHpo
w+8IwC/peMB1llAclpvy6GRefR1QA6KUT1Kuhum7HkuIC+AZq0LGMsGq4d//u/JtiwK55QzOPP4+
/dhXgeB3ZuQyO1lElxAlt65J8EWtQ53wJJLERuGKVcCBocQ6WJTWHyMOrnSwsSupQZnIAfNuk9Oh
cQV33Ma8nGgyBCD5TBX8ZnN+MX35X3+IH4ksNkjyrLlz4aeMlIHoT5sn/r+DZ9I4e4yrwqiNDfQD
RjOtICZWTnjhlr0ZSryT5YANWWp1l/P6CPmv40BdrLXkFtW9EwdvUW8h+NwDeXCnimD8xVkVsONv
r7eyvittPIRoyhSCTPstu6lN31PzfLqx2saDfJLK1Jfspjvc+m22cOmhBegMANPVP8g98H+rtG99
1TEhlp6wyXHHRASa0UhwbhCshf1Zt609MMaj3cpd+jTrmhtxdd7vakq2S96fKDRrv9fSW7zjdxvh
SIxMs4ymHsurdNVH147avSrNrQoK7QPPHG/ZHyCGwIwufEYV+P2D1fnQcX4E/i6REmO2NV+O1xT4
EwLP5H4tTI/8xJu6huepleq2FN9L3fTDG0PoHm/iL36XQsTMPWtjH+BxBOCuBZyZBnbL/5crGHhb
KGca4Uyc3EYKMgamQzE3CFzBc1pHeXt7sTscaVDzEn8wuu+N/5NeoutiuN+RM2zT6Y7BiFSfPQZE
3HkfsSIz/7Vz8Mglu2I+2w0YPrbiwrSbBspLyl2WLUAT1R/Tcfph1QBTrKLF+PEphQeJEutSu3fx
ca7JW7/zJch4hh3ISwqi0ub5xnvWHX0WaY+HzwXRvZGT+LIJMlyQ5wTiEVjEm40JP7fD2m0PAujk
DkP8jfT0C0m3ZHO99m3sgrHEcg5YKlxHErKjMdgnRVEmStWZGVis5XcqKtxxTj+Q8Wbz4/4ZsCVN
aRjpiUDEPfZel+mpRSYxkSLMoyYucysTjn3sECqSn0obBoJmcWm7nD/mEPijvQNcoHiAUHGUyhgY
uWVNN/J2v28mvWZ5ghTXjaYN/IKgoLUP5Ag4Hp2EcHvR1bbmrF2AmfesrI8BUD7ci37ymzEG82Ak
v25+VECt0FVmiZ0fSu0C/woYH+Eg1hf2611jGO8+oKPZRjkIgpyFB6Bkg59YW7DgfHx8qJcJNTYm
ed+mu0AYMy5Ez8mp6/fu1u4bhdYkObBKLQIQTxAvCVcvQm9Zj8M13fUVhlB0Ugf2nmBKs/+F8Uv5
8qOxS6H/1+v/eso6AV9FEnxrau3mOtRTHRhQJXeS5v/4OO3COJ8P7c/i2UI/j3TE/jVUTB0Ztt6e
RaxkwC2I5JNBmulRzhW1trhsgVq0ZTvLb35o0SLX5jnCVWw8dwUXtjBc3CRwwpHWDUtbld3AF8+o
/jU7SMjB+lH4hEwdjNUohR64sle7vaDFuo9IP63/xtIsteIsHZ8AO78OEUNVe9Hvag5jwx52snuM
KgaBiFdzbLu8W0tT4p+XqzFGKf3staidOHHNEIVRhGhmvPlFVinMZz9ABwV3gPJdM+LGgDUXT7kS
ZgFRcOF5VvclkotogzM3TgDcbNlQUjGPzwbok92KQJ37UjdrTpGwroMhyXtSdKFVMrFwQvkqQUX6
NKVwcxyGnJ+xLjgdHT6eAmMG6Zjcm3AO+C+A1cRfxFvTe5NU1kJ7E3RzpO0vVXFnnZ1LWgTWZxhz
j2lpi1jHrS2UmSSUOIh9U6k7/vWpgF8AmKKsq6actA8QsMvBQpbUXWrPNJ5DYzuNSTI7ReM8PDCg
KHUGdYxpPeju5UDijShuQrhqy8UtLRwQj32GJFw6dv8E3MDXH6O0vSE7GnIe2g4YUKd36+4W11ZA
UMkbruPTgFlizOO89qYXM3GKpeLK5LAnc/zjjZ5X6VDzhbFb5IAvOYY9m7f8yf/KIXFZ5193gSTQ
ThShwr3jg3DQCpMdAB1UleVi+NtujmNFvqzEmqrx+EEkPvEIL6D4GslIQAItzXDZXnnILVsgf183
MVI2IKowWaXt461RP2zObfnwSRUO0vwyajGoMW9hZbwJIAjp0ZxMnMuMrNX5dlZVTBJW21HSDnmz
EDzmhBOjhKRBAROEH13oHRC5S2Gy5GFVsskATWs82R0oHgcfk9iu090FghOcBPvHD/s2Ox/N8jnv
mwZ4n8xNFsau/QCff6hd4DOHV3MNRwYiY/VIJAKJF4VOi9GT1o9CsS/LF72Bv6SzVCSIKNQ6B83n
5Ae0Vjg4Yp9po7ZRoEDIia0Xkk+k2J37zcx6mVWx8HonRMMbLr62MMZpQ4x5HaRjbg67PaNK7eZ8
vu0MfWIQLa+Gwv1UUvuT9wutNxYv9M8TP4T81/3k8Xv6fTQtBA1gZHdj/A7sFVUGcb9V7ottDhPy
90gBch5InMO0Gc3jVw6D5UkI0vMkH8Fz+ie3TR+eQkK9XGuVlGijFCxdLJuT3mUGwEGjJCoDCpk/
nZdB97aU5cMRHc8Zz3ReHV8beJonbGx6atETIbuGJ/AT7SKaLsJwCHMvohM7c7fR7UcDmIflyX7q
0LI2jgx1FOcMy9+7/di85NpVtwjkyetbAkSAUVrdPZ8rH5UcVqE/7FeS0qOAfnDDxLExxDY28ICz
nASA3JkSIPaHOoLmhhAWYpM9QXnpwg6r6v8a7cdecCHP/pqeSRx+BC/HPH3U1Hi3btkgl1vJZ0a2
8rDJx+d/qUpr0HJmuEFsyH9KJhwN4iRq9UilnjslGSiZ6ve1ZKrndaUFfI2LABaVaXiCOYc2xZNV
KLL+GqyPOVrSBZSZIgJ/kR1zZCpf6228rmXX9B+km6ZQ6pUnsekR/JXqXhlPHGx/kj7v44+G4HPh
zgodGeXZGUG6hjb845JmnG5vAV6UqG8jLc7k0Yru2YJo3K9oo7HV5axtM270FiSw72mI+6yEt5JZ
HO5mySsFOwB2JW8HcoCp9h034oO3trwKz2pqovnysKRJn6i/dAW3eJRhRLAkoPgah9fJcnLoRqF9
upNkkxXZ362JRpgee3GicWqVF1WaXhDQ5esRG6f609PvFJs2YRQDqtTKK3nzXvykMYjvkJYdxGIR
wCo0UKpNsrSTgjEx7SzXiDrnjvy4wRWgn6b3KcKligTY73pyJpScZWyx3Ox8bCInZ1tDKNg7j1mE
+ofZANxH52YSNxo1ddJzDxAkYbWokvdOqI1C4o5EkjZoy6r5h7qEBPqP2WQoOW6xV/ozPGgANIfk
lvjPvXfLm1FRYeUmDQdUX0/48wiP0mf5aHKIzN7xpq/ws3n3s69kSXEJdpQG2u98kL5m6OAi5HpN
OJUzH2Z+7HupdE6LVzMqnIzCyLaO2KkM2GF+ax/yXYS/4sOLu0XFSGirrrC4i62PDJJS214iVXap
4iEtAcAEhuAwUi18nWZgR1a27bndSn3Jy3OtG3Jn/F6y8tH+E+RAS1evs6Bx+ckWkS3ilNWqIs1K
CgXQqBDR57LL/j0gOqvJE374LtCWgH1loaJLZy9sDyNOfbb2TR+EdCKpBFvjlDpKv6fvcYkClURS
8OiQHb0oYUdPyCrz/N7mEe7svONKMwylyi00AflbQ9QlJL95ntsjDH0xlUC5/k37FHUCOjHkt8pM
giVLxmoyAu/8GyOibqkH6tfOmhbwB0kNOUZXS47bHBVmiZly4CVIRQ/mue9JMiPY868u5BzIfarm
jBlUOK8N3FQMnewLjQ5FTYsGsyUhCuN3HK5WCan882rSMDr70J+KlATgxuwwWNNuS6xolU6ajFi1
K+7V9ixHyx4+zxZzQM7mCBZVctXNhsDirK3hRkEH/PNlNDzSFFfKAV2HgMiuH0gsBEAfpBNdRDae
TGjczbuh94r7ArUAvzhaaahWDk1TywjN9wnCVpg/OBICq84eC1FpI0NHxhEvTmpwNDXY/b1S+t/m
TfTcNz1FvUnoXMV6apoIXnfBrFVVDHsGymGIniqkH4kw6dFH+gDyYEVn7pJxlCom10idd4CZktln
I28qoakeyUAwVfrgeiAinHs05L7DkJlj8a0zyB42ORbzDZnZ0cKSILn6z25zseSfsGtJydY2usKQ
BLBWS20ZdwJcIyBgAVxcxR2tTt4/ZSRpJ7AQIyrcxSTMgT+R/LLfkSzCbNwFv2WJ6SYmIKozw3kn
sn9omXIr7OBGrIOJTcqIAoB6ZZ5c7hSqSpBMzZ2X7zVJ8NLPbUoqxf3zx4Xf/d4l4ihPPNUzLCWL
ZtpS7lLcizg/w4W9o1cWkHN1ZfdbfQk5UHZXtgIAP+tfZ+OW/Ld/qQwqjpY53toVOringcElRAuF
OZ3DUgzxz87AMr7Oa55wRz9bA6/Qu8DDegDDB+wpYZSL12TIgfRRfqkGmEgNYu2zL3bjSMXd7EXk
iramiqNHFhzYwnp/qCi6sCdt1MZsM2gqLB9zXL4d3OV6YtustVsYuv10JAkj3I5WVn+aQP5qYNak
Gd52xBS7Rqk4tcEcgKqcM2OIsKmGYSjaYuiUAS7RDYqWoqZrt7rzDsrQefumgzs7ESzDzGzUXC+d
V3otCqsS7BsZO0u7zKvrm+aAFO9AdK4dFDPjKjTRO1O1J+IV53Seksw7GSzbLU8LwpZ1ihFSEzt5
g8lTX5QFHQspqw5B3k4rFE/x7RjtD2HRVGgSETeHZnpJKhs3VqIm5ltgEuVYMJkOtU9Emr7NTZrG
F9wnsmV75gcsexIelQqH7KPLR/ghvvOQ5CvKbEteelxxjUkAPC6tj50JlRL5iag6KcE/Z1XS/Gw1
kJ2OihqVPUVXOFjDq86BAUAJfs/Be+Fr14HPgjXfXuDWdWa+kloQeye/Oc4RU3sbeGOfsmDib/BS
u26/Sv+3vA2yeMYm+Qx0I/SsmkkvHjJOrDw1qZkF86jKsbvgjdFfnZ4JAh+MOy5NS7tb4XPdCN/z
ieGHmdIRNPYSz/aN20LxCh9casmKPR/iIvtiitH0L4SZjr/fgBPO9HS95IqurFMF/5bRjpk8oH1K
BZCYorg+8mIkxhb1qvMfEaeWPaQFpoDA4AZHy/sbv/YbWVM/zZ6fjjg4LH4xR186IarfFP0/PGDJ
bjLO0Bl02HJJRRQggJ+5ueDN4ZFnDrvCiRaepX/Y1bDknOqMumuZliHhIyRu4HUSOOB9qT3Lz+oe
4OR49QzKWJsC6y2VQEu9k1Ha5+7w6o1MjwsfEVvbWZOaf6KpHPfKKGK4LC1qvkZ8kf+jJ6GKLl7O
dleHs6uAj0+0JiMM7j5RsAccX8L1pmatfr1lgRwAmkvk67dHorV+ot4D0tW7F4tqxtQa5Znf+qWN
Ngmo5i05nR4t2JvdYQukFKt/YGQ4yQuK/NLQ4MPSFsLOOfBMg0gAbIMth3MmehG9ZByMdbDozEsJ
yAphDuGDxzGN9dVi+V9LppCfTWpDfQzMH6upo7hhttQvoXk2AOfiUE++WNEBapg2jf7iZQC8BVAr
LfpPsRqxinZBq5Kw+9obX/y93Spl1L0FBbYauR4OIpR1xXcZ+hQfr7G9d9Znxj4tJnGyFKaJZ8+j
MDfkdHxiRaHtGuGILsJVZyLSZlIRzgyj0QcTFOWH1F8mFXba/FIGDJWldSIKYlmT2YKgEVoPhnKz
uK8/NVCFUjJyop8wqVWTyLn/ZW3f5cktsVyUJvRtY5ONbKfT5+NoLV4fLGmVmn1Ij2KwKsUHP3tz
rVOqGtFC8ln826BldwfkQu5wKkPzeWjyBILPRG0yXnJnMZtvTHXm0WaAuRthop/wx8QapQelIYXF
VjCA98EEdKlzEhXSo2i5M1cgaBE8bSmslu7SFdlxvgObOfUmA8zmBxmha2KoAdPIR4BNULgnRVdE
+F+sIvcszB/LiRt3ZcBMLvsIyug0wiG7hdu0hi7eG3S3chgBWCc/mFIY8Pgy0NltPb1iYZV8HBde
A3pTUdd/eyVg+C0H9p4w4nIXq30PiP4pS1kcvMf+R/Zv62+IWRhqH5baIBIzFkmJTp4A99yMaOrm
xHAsJd22uKN+USWKG85zYHUEJEfthc8vJLSKng8qqqcBUcHj9hC3ut0FH4zoqXOd66e4NnjWLSLM
bP1/aRkZJOLgfkbR39H0afEfW+Um8fecDnHt5nOC2BoC9HK4hCgRSppczy5Z4OVj2IAEXf1D+sLH
EQldjrzJ46g/c2J/576E1yZKTwTNdWmnYFbNKwTVXA+vfw1GSAzfdbaBTwlg3V5Tz4PLJynJJ/VR
h6ixbAq3nNSlDjytOQduGNsTyzq9gig7vkkJea8tubGGh59Oy2XOUjbWnqMFCIkDB1s/PtcLmTTj
0sQorfwllrzp64OEh6fViHQlj+QvGfJJ4HpsdCDelZM9KOVfXIReB3ZzUzSZFxqAF8IUliv+L+eQ
LWlpavLqubPNgBaSFam8WnGN24G/m/F2Ho9qnMZEkHn+jZE8bOWe1hrqhzmVIRorRrMkmDfYYoAd
Uj7lWrW4z/OpjX4a9J3EldhTbuV11kJucxw4JgQI/BUkh5NPW6kLiFMVJWbh1qtCCn2YKp8Mb3mI
Isjirqq6JY09WCWdJ1mQ9ohQqSXjLTXtWtNDO0b10H3JRnE0yWCoN05z4qwMStXBecsppfGeMTfc
2tNHCCHgytlEmJMZMFBsKUN6e9Xnh+mUJAF1ib5Tn7LNxQJ2H4ZO1OzQC6E88lexjd5ARoVdJvA5
/KpCHfS39u56+NHbo/XaU6/OZNfgj8ACRMbhtAURdf9mGHG7eeIlTbaRkHyhMPnL2A6PARvWyQxu
s4M3LOV0E4OJjcfKzYZpm1jRmVwRWaZrb1+93LD3sGAZxpr0CpBhhujm6YH/bnEttgeCkbvzPV+4
j+GOtHMVqjYGayxRHCV/kxgl+INHhF17xUurRNXu0cr6dYFMW3P3KXRi94jAKKlLBBH+z+z9M7V2
u9MBNN8nSMNa4EWTjjtSBXQNamUVmH+bY2zUL3ubXepo7+pWSU8YAEl4UtHlQyDPb/Zf4LhLsR/E
Cj+hBrNCEa/MpSHyrghTgnFdrOSjye1VRzEU4bXCg1cvhd9W1YtJcIyAERV75PpI7RA7fK8FCpkR
0RrNM8w1VHsAt791AdTAnx4onLlu+Pk9EHGsrMwTi8xxfwsMBZbaFs37VoM+2fXkSg4ENASbbs65
V4xlVKeNiAKk4y5FbT9/EbrdaavaqS53DCbVcmGfdFZ8UQcImoxYghrozGZ7zTTTDl9AEwEE9Fwv
Dh+kDi3QjDsn/tE9z9zsnysha9UKy0R8gM6qeHHZ61m6c1Pqmv3UCWZEKyqXW3ue4qbZyYsXAx8f
6fNZgjzzM3PaXyzuP8AwNItwZ/qB3mQnuxIM/AVBJ5Vh4hjPF8dQD6RoMvUgYBHeIJzZrtbHx6is
o70bv9+zApTEyn10wnTqIg6Ue7MmtZvq+oZJMcOVMsDtpAHLi4hJenc2w6tjWOq71ZQUkmqHSMG9
fE5wQ7ziLjaUbr4Q5eD6JRPaXRfbq25LjnwZkVCNCMW1iEDIinjpXyajpoczySHdYdBs54UXYrrN
+k/ALk4ReTgkbbBCPi5OjXDgL2xC/b+djMRAQJRtqQBbD3DZqcxrJBJItlnFPc0DhXB5jGj9pgqT
n+LPWcro/MSpPkq/gA6gEcQta8KAuvr84utEbIjw3YlY3Zs5E39ZBYEzpgcB/y+h16C0sLmW8qL8
0Q6Vdsniy5qbADHDKrVv2yJ4uvgm0Qeo/AY+2WzL0u5pC/0gpVsDrAF4/7TlIBovXpUM7h0TYDhg
76e4F8B2URyVcyjdroEv6TQrKmkQlCkke2LnnSN48gt0wylgxOqRzbzacVVeHMhMbwcxUl4J/RGD
ZdP01psp+cyaUpARL89va5bS/f2OX6ZowscrZQ2UCKfFsTXGaMC61x8gxdrYWTJ+0xIHLcm3MjKD
5CYoKr/7PKgoXkWKFGJEMwBlly5vREpejtbHoBnFbvFcwHmHjG5JuTQdwW8DFMjXO0kLn0XZrgBe
Fc1tN+17GQ42XsHBRdMC2phV0f9PqJxgSoDl8CCyEiylW1U5nQk1uAJXc4OaHLKAhSIhtMCcDFmD
B3yRZ12v+Iz/Sz2827FEmV2wPat+GTKAnIxnSJNhYeYn4V+q0B5jggs8JiP8lKMurutbPCD7IhaA
krSXv1zDJSBsJsHm4evRnGewsf0kFRMCfoclhfT060JHtDwkKG7CBWa/I0QV3BtT+TjsX2eVHRL4
F7RF7qrqGrJa1B8aR55k+pAV+r5HrKuzQKSfqEpQ9mbymTXpCuyJOUVd+R8C46EATviocjsDqGZf
0KhT+sO9gO64DU0WInsVOTf8yX61hnwR42NjZsc15uKwugf/DPu8x0mh2GmfG70fvSL2wyC7odJY
cwWJ206R3/bs04/RDo7Kfda6DKJh6B3HvJk91ec/pLkcPshG4ByaCkg6Nf7PvR3dmsUx/fLCRWfg
u/Um1QhFEMfX9qbpTz5JQCYeyr8zhxGDDrDvFO0pMxw9fJpzy2kp2l4SPt89nMJ1SurST2URvMvH
dhkeGLcG0MlttwCM6QXSg+AKBprY5KUJhXl6iJXB79SB0TARQbsS1t8V8dQ9rRpQzA1/wFAuICBF
CVH1OIAxf3Iv9OEK6pNglnaLm4aQOVlpQ9m4cT0TgaQmayd03rsw51us0k1iuju0ap5M3CUaMHTg
R2NU2YA8xyHhlQ9WhFWGKxw6lLgjU96SI2itSLIv1JTzzyHvL1uBThOVnjCSUxkqviXEtRspNs5o
cxRTGBL7ADNDWqldQUe/kp6maTPvwRDD+HPD9COw18GR5hwBuSMDySE2eKMod9msIpKGkdAdYjW7
msuPwGALRxqNStose1en9k+s9tMA5ACmIZQtHXZw1PqRxhkr++nQGXx0AVakNDXVOsjHy6P/+PWn
lIO9+b8D5n7StXiD0gZVfwq+u8PVG5Wf6skHXuSAZVARkMcbOPJPcun7cm3ojBStaFZuCCFw+C84
KKajsgA/RvH9MuUgbQ9qF0vWQAjMjXuI+bK8G2+OgLkrmhjYCFF58eAzyO9hB359saLOYigfYwtM
90d2Q+TEzXAPqnyroPz0CEeT2LN4xIP1C32EJm3eARXAJMyRwg7MqweArQZwazuVPHOcO+BFQwPq
fkSNQmS4ZLi2GDhGzZrabBc8kDwmw2RIDI7/BcZwpGU35r2rJQBJhI+29WFkur1pLbFfbnq20l4B
g6vj0rxZACa0CjXjRpYceXQXZSoX2u6YEfSgBL0Q9vvDCMZFQZmZHL2pBXggKFleqTM1ypTJgtGO
Nmh0/ApbrCwJ1zdB+wHXapjv6Jro/qRdV1pxUBVcM81SV8O7HznEPqOswfgqdt8nee0FIy73BJEY
2ARjwFROCkT7VV8ysrIdiSooqEzmqD6gj+6PK+dv2gruraVyBS5vihNDPVuMP7ZerbJkcinn5VTJ
k///hXexM/cAwYtB78QiVgRSqYbJ3u46qL/v/VNaEvJl1cJHEvEgjnmZNfeUjVcJY5kU7D9uInKV
wspfZaq1t3g75T5NRs/hnIOw84DHeE1e0JETsQo+sja7WMZrTsS7if/+zQk/HvWoRaTIZ6w5JCLH
N+PIiaExr3BV2a45WZYyAmS4IOOqHzET6gexJN5GuIDoqH1glmDdFvJLuZGnweoMIL4fTzTXD15m
qZbG7iqk4H2BtF1sKiiC+KvUZuVoR78jgFd34DfTvy0SxiLTdJKwH1Yj4s3ERbC2k/VtR108AvAv
Npy3NlNxdpjGbs67jnrj9EiRliX6dyrFvm6K+hibUdSfUlOxpQZgOQE8yx0pXu33ktYOpBoOBnZO
V5mxDCsfMMGFb64kJuj2FBYrS5mBERX5CswaV1vxZOsuO+7KMyxmBkjaNL9O6ysKqBb6LpfvaVou
cfJifKdwjWLRHd+O5WOhYpyX/EWDetFHJVXNkJM03gt4tPDBN2ApRG1zfmv3XKo+fGvxfYTkAN7h
uCjwLx116svZ0M4a7hA1ZDgCqMMybxhXrRnHsVm4GQ+61QKCtlZ7aJBw3cTYVu19azIzqVXR0XHM
cdOILd1fgZanjP33fjPsMyutj6ty5z4hKzCAYSn64OMiJg1u9j+YQraMkK6E6N273IdD78MjJc0P
7x3fPKVyOaPhWWvAsIR2KYl6rukspir/9PLdQFgoLtIPA6LSZG23g7ZOTGX8dMChwccU8DVyE1RP
gTLXqfcVZrmHBFn2pE+o+VL65lFU2DRefB336s8uGgV6CFjFiblGjN88hK7Ix8wrq/tguosREW8f
UsaFAIYXzeNN6jeOTT+HoZSVOlSK0WbNHIJ3LP6ie/6rLWBR/fLaJX1/60HtEXCY4LBZuAzN6RTH
5AHaILW7xrYxQer5GaIIot9tCOx8z5VbsWbjSpQ1APF7O9eqPQlz++ef5tNsVSRovGMmOZ/x8Ki/
NklQvcc0BYOruX+Yehqbho70zv2i72L+iFPKCedd0uRIMXCjF63AVm3FfXmJYJIGLMS9dDmUqQDc
msqCOhKK8InUsXHgyFMQLHHjGCopxAPaqYVIApxiBjR9IvHIvavoigDpAwPMn40wfM4k2VJ/pY4b
vy0d2ZL4Wu7WJnhi2Pwl6ex8b9JYi6+ALaCuRJbhDYMsQTgcJ5q9BOvIxAf62pkiB1HG9WWNMQFW
yR+ednfB6q5ZDsP/Z0E5+CMqjMF+6trrjdUz3Tqh02bWQ3j0wEAkXz9Su2AwZgCqC3Z+Iytr10G4
SUYXnRzYcDoOm6xfGNPzbo2S5mEGf3RlscHViC/7UB7gCH0pv5aZQZVl5LwGs9i6ChKbUTRAZmqp
sxBC8h+mbKasteky910fEpV/MCFbztfSKg/UmORr0WpK3Nuw8VcSf+PyDiDsOZ902y+RyDBpAQNQ
xjJLfzx0R9o5t50ityfiDMiO9bnv8tYYT59tyr0AoxTVtEILN9JGBvXXw99uvdmo63o7T29M4nR5
hswYLT4RJP1UfXKSU971MlnXFO2Wxl8tIShaMESlezqPoYpDT8+6Qan7ZzU6Z58qi3Tg/dvEM7SY
9JDbu0/FRbNPpIn/WaS9gTHiV19r8M0cSlddJoCJz1TNFyXYXQT1dxEG1BBZ3sX2YUdYD0Z7cHbq
JbCJeESOi5/dN/fbdRZBz2vghN6Eb1MWF3YfmuYgTKUPcbiWtm2yV5uIPIHdFT75a9gQfnlH0xLV
MZyDH6QYFJ5tOHduWg5AEhjdUn5s2el6M6nBq+tjh8IUpDf8IcXrt/BjCRvknnr2njLXA4y20Mjg
pjqAdzNf9jGQP0Zt8s3RdgR9GW/bk6xi5MkP0Rr0TpLRJW7CcGudVrK9So9Padrusqs83o9Ye3bE
d0OEDLLSvnc9NHA9bwFg45ZBVJXUZ5pJV5DWuyjn8FtNmPfQd3TeFu+CU8BV+DOwYjopERdBuXbN
vMla3GM8Xoi6eBjmj+fuMx+eraeSL5YGtlQMmVdQPNOPvE4CXEhZRF/QVLUGRYSI8twlAY+vVRTu
+PlPgDfii/4Rfc9T/jgOjKNbwAoj3Eq9M2uv7B6DbpyV2NGD2KO02v50f6+yLToZvQ21MPAWiXLJ
ZxElUtPP7sO95vDmRIPHeQjrTSzu+gCPtFpBxDV5AQWCQYRIVjB7Om5bdRh1O8dmirZy4Y3BFoDj
BcC+S60D2pK2URsSKDnpdt3Qyg/q3Cr6O5UIMZWpQNjofuulGL+//M5CWkBnpcmEeSyDJngsxr0L
0tB5NhpF/VLzI2MpHVezF9Vt7qJtAT9tKxWTdHhWXOAAcOQpuCOkbibp+aMRpnDlOQn+3b7UuFD2
F72yaGyucl2KETkhsSEPUdHH8XLUlWZp3THFmbEX46+kZlTwsY8SO7P6uxmch/PXDmNLzfCwnnfA
qI0e2TfM0os888oH484qY1px93etRcvb/65nkErGD3G/vOZ8qCGGWK0+e5lGP0JRDKcX2I53bkoc
MEu6enlZxzdJtybgRQkLDU6EdqWmvLgXmMQwpe8re8GC6VFe1FemSp76o/37r/ekiQeqZWB56oSS
V0KpBD1ff3nR81Ryzzp2T4i4HNBo+NKgfoieJr5XDf0OKdaM51WHVJiCHKuSCFfAS3udDT2lpNR2
bYTbl6xDupD6DPtQTndsy0ZsKaLCxDABvuKgrlC5rm6To1lsy6I157MJMzkJOc5liITPSBH46Ges
uYPk21mVIacVSj+jcBntE8ws6cPhBKKhoxImQHSZMOOU1dGqIASXEL+/UJOJep3QQ/Njv1Zv23Mz
jWWlpyNKv1ysenmpMf2vOo6XrmM//3kdMrypYwxh1AtElO8pxROlfZEC5eqOOCKT+nS6FjoAIrnd
S3QA70fo8BYNR5bSkkxUBSxvQEUDfZssAAYcG8KqjGLm+Cr+qpSIf3zbhVkNltmBdyPdCbd+pfDa
VYmgYFXh/TJGLf7z9QGCdwsI3NQBGUJGTt/FYJaGKYS2u0IlJ1BOoitwoDmgSJnX8blzaxOy/njF
E5E5U28gbzdjwD5FJR16FAmZuvk4gkUFmWoC6IdIpe7HK1UYd1733cZWxHgw+ty9edUKk3bFtW20
bcmzzL1Y8SdMoUnnFP5nkbty5i3RY+r8o2O4nVc682L/1jV0RdWeBlicH3AWTLmUn8iIkO3m6QSp
IoCIHi7yKeYLj46UuD1GI4Qqvd60XF4jC3fTpRV1nSh72t5Esj3/EKmMwRRpcxBV/6/vLmyWBKwu
LgxF97/bFrTzeqBDRU+ZlOFuQIOS3eE1DranVaZ/waFP2ImMT96PWJz9Nowc+1D8/uacmyuzQv47
U/mY84yl17M9NFD+sEGeZrdUnsuJsDdo+Xfvh+b/lCneYapgb3SssIntOJlkXVmhI1hIpeCTqVHJ
lS+f/H1GN7YNtoHt/sUkr4DAQWbXG0mw/rERY9UdIhjULEgUdJmEF7YICU4lVvuREnLcHhVfb5Hk
GB+ggZpta1bckfYvZhR+mEHTy3BXlOmwYcjB2xoVmoOQauaawUZ/Oa2H5HHCKDMY3CFi9JL93RYj
vc9cbW2TmUj2L+k4fmH1ikmPzcZVVF2OAD/wYuucjJJunSPtOOxsrC4NijUKQXdN4pLJ1b+YTeaJ
uTo/bQ+kW30RVTQbcPF4qjPnoOZU03y7FYMnmykUvyumM1LRhag4OFqMhabX7aEon70qVUBXy8k9
pFbhtYwxcndvL0iSpBAnkYC5Q8nj/32FTe4wIqc5iw3OU5rb8IjObrKKJHPdbLl1j1N/sIkOHRWP
UNUM4Dx2tTjR798XNBtoTlkEtdptHE/R0lALwixD/F3sIMaQ6znleQUHzSz0v9hh+fjgIWLQClQK
T4opU2mcULQvCE44SI4qbI1U7lu5yG78+oAc1dt9amsXNhpuXCxPmRm3UyLt0+yK531tAC80V3R1
txQaC/Nx2cX5jc3D35BsIhV6M02+4ni2CE1SMSYZKjV+iJthTJRgYzduFWhLdXmh/9HsxgEbbZgj
HSAuVrXzalFnTGDyEH3lz+xV1fu+MkTMYn2ocH4xafBkYnv4r99OmVDChxnSFo1f1XAC4ROv2Kuy
VfCWu9LXsWu9ro6dXipDzvF1MnnMJnpUQkK2aypVWfhv2Y1PNdeVioEkJNmEsE9hLOn8bkzqPI8x
IELTeZwuENwFxkUN0nEiOpT7eRY0Ne3/KQ2JhNDJYdMHPTohH41K1t4RxYoybNoJAzZmfeg6CPb/
hEOKiDdc1UhoVoU4ou0WILt5+4zF7fY8A7eqR3rM307MCJZtnSiPGQ51UFGYvXRPDIh1QG+fkgun
GS8yFBVUi+yJlOuKbHhwk5er1mwoCphUesU/XiBhOq0KiKiHJHTa3Y25q9fb1FB3qa8u6z4sBs/k
qeg44KaGl/3IMFFPt4C3WI/+LmRBLhVxoebLdtX/dY4ObJ7eDrBfAS/vPhbARfu8xiLIX/94icV/
qsDLmyGYli1V6OKyYz/z/CURtHhwCkkCd7CnQCPbmBiLmjVGCDHPX2QtUApBiHcZlfF7b7ReI9HR
G+lGdzFZjHIZLpMzLYzNaVgcjHIItetBcKKvUqPO0pOZtYHeyhlHPQdzRGvqW4vwsIzMGzGoFY5S
laLsGVb7n4SzXIJMRTUyNPPrJAMYopR/MBt0c+HoyVaYWSSOs7LjA5wBZ15i1DncguLBYmM4g++B
/5MoB+++ahxy9n2nkcC4yjrE3/et0NpCsdpKjfKdpEj95ZD8mtBf2lHLg1ZMKCp0Mf8gvmyfmKd0
1xjIRcVig37GfXLBnPFNTMUw5yhN9DKFv8OZWy5CwDNE/4KSMwqR7Y8cyZs/abE1fU1tq2gtS2C/
Pbp5kGI3SVOOmGDfL+Eqmh5cBXousq43/zf/lEcKKisu/R9jiF2JAlGHvg5s5tqYl0SEjHj+oZWL
4HAmTvHxpLkdqdDAXlf4zkQUZT2tV/GBr8HdkfsWdTo1wR7eL/EiGqevzi2WBJz3+r+NcUmJgOVV
e34rcAmVh3KxltGgUO7Xm+YbG/eyL46WyoVSJ51fiNY8UoCKV9eCkTTKyZTTuzr/P9NozXWr1AsZ
qm9PYu0JGW/IjrSVSzcGvnZ2kG4vA68BZNBZRF9okQcwzzc2ald2/WZwiMYMLxO8em+UKkmhkUoS
WZPBigzJhb3FdYb+km9zpEA+FomteTpw0OFvejMi39TKlfXGjg1z2LyToAnDBy5yZhRvwb/zgWmo
pThYNj46qolwS8/QEFIRpii0XdJnTxw6OFzxgiuQIAwJ6ndz9u+xqHrl81Z0KxHBOIHGQweZYl9v
hpw/aMNXk9RVlpXCMXaX3VDvUFGAQz8VmlbPjqtY6I10b/+SYEI3EuBUq/OTZwxztnP936ndirj/
4ugQ9kdOH5BczfEL4IOkykwnSAy/ijxD4r3z0Hs/SfuAShlB6VBqZKPR1ZlVFUz3TRPx7Da3w0iw
h9O0LbNdYGVx8D3DHoQwDhlD/pcwvFmZLQklHGiV3DbgXudP/yMcc1H5GUwZZtvPH9zV33NYmVCT
kYQI/wtcroL/ASNU11baNDz02HKOQi3IstfaznUp2UJE7D3EBXhfLDxHYpjD8Dam/1E1R2AHcekE
HUDth7Sak4ih6292mKJjnqOt+WPGlMqGibbFTcdU/zZnaybq1UDkRltWgZScKtX6DU8nBJq8UlZW
vcNKutjuBgDAeIs6k1vurMLbXO/Wfsnpw4gjsI1/7197SbMfIz1XjbJv8pJ2c2VDqYUFdEeC6FYo
TxNZSxhZscVEPBtB0b8nzu+0Dg34pRAUq7JvUfw8r9M1ODHJCBg7WHU76kEHCij5QIIX6E3/1H4+
SWPdZoebI4pj4LygG8FXtuuq37LqJHIwrIlyCtc1A+Z6rMmc/xZy9L/hKZ+54h2zQjYfRGEW/HyU
cMdpZtwP+OlQRsT3RtJJ/NyB+wMx8PyJiGWWz401N96v0d5+lzG2/8J2R80ZnBQicGRqpJOg402D
GLjr9ZZ3hH9uXJRKrhVNZEmLxBUuy3kxENUUTBq5vkXSfQVzU9J7JJVW+/OC9kM6On7eAs1Egqgt
NiCPxKrchmNF3Yp6GWzs5wIiWHRpv/wyPkrBL0HFpunHo10loQaQvmdknwbZJlf2x4WfTpZJDVVb
XOa2zRMxl0lKT+joqQFqEJGRCeWDs+uV8lNGkJuKK6l9GJWQzKHJPWfD6tHB7bGsqvrRDwAzZFGv
3mbV6LuqbidG4qc9Lg1x15kamCMWmjT1RrfZ/s8QSYzReZmRnUVbJPaEa1TYTOpQtDQYhzJ36xxy
LeUcXeeExpkBKAK9ScRU9NoHa0HnJNQplsKKoZWV0tzLgQNxi0dzNs12/H8nhZPT8xVnT+guWngT
D3MPavhn5R65eydsAsGlrPncF15zRgsBHmk+Ci8FSnLHyr/gP97uuklo1DgXnkhO5VEw2vfhkJ+x
vSk/YC88FLCk+K2KztNC+LVig2sgJQAJfEVQ9eg6xE6u4/nctkoFP1k5MbCCQyDFY5PKKlgzsbg1
ovvTum8CtSD/Rna3Bc333F5hPSVdmad/EhXDbbSxO3TKLI8kThEUCXDkWE3XeKkjpRwT3WgG3zF8
J57aOqe/3Ge4fdDscmoiRd7cwYaiasnynNWK1mdeqfkSoFEccJZGAzxAWKB0P26rPZmIhdEpHhq6
wR0GKsDeGpXdaLOxJ/9aMASpVQJyObeAAFuG4wETnBSr4NzFZyiYc9ZqxQJY+usA2gPcYT0RGBEn
B2eSEj/K2pXLYAozBjzAugoCI0uMnzWpt9Y3L4jLTgZ8wFebSrvwBQ9B5e4g20gKl+0f6mHederP
hzxONa1OFRgHv5Q/6+WUiCOTo11Jbm9rNCnAvOhkdRZI+yRLVWC/6wAbJZQjtJOPsCse0cCm6IKQ
qXquFQO/MPULVD2foMUyzmRCIChHCGlGecp5yQFFaVAjgyZCHBoHhR+Sss+EMggYv5Fz0xGyy0ws
pUaUAUG3UcfteBtynbP9dV6kkhftXgklqh7+f+aGpLasJLSclbcmXu0Xt8CY6pdXkQ2eyNXWrNFQ
coMfjXslGf89Oq5Xiz2B4R2KVt+/XfFGbvzRlSm//3D8D52uGRo3aaCTzQDCvpLuemK3Oc0HEV8d
h4kqLcw/yyYgrMmSYmPeaM51s4PKZrCmpvN02oGFcOXwZx1YSYPonF1jXfLH8wgBiNa6IHAE25QD
BM0Uz6oRblB6KJx5ufthe3xxsZMb3q0kNvEIUAo0fuA0Az8PKs0MnklP1T7QQWsJmrG4unPcWJL0
p21x8r7Tveur9FOQY7CP2uYJaYUWghhdY9wvHeCRWaqsfbIGYXML2/doOW/S/n0pnnTps2JjvmM4
DMusaoA258B84U+2C3+J4Z5Rn7D4Rh2B2ZP+FC5rt28wgUjWdrNoxKkJgXld4TxHnLCkDRSj3eg8
XtzG9fPQQaSYyPdYZvyKH5LiYT3rnAZKVC7UEqOpRZ9jnVGP99+vGjh+2qRzB74YJD3d7lfFpMy2
eCmGLhOJ6d6KqQExGIQzBOgujOdEOgvw7aSsH0qHievAOosIeLiT4QQrSJEg82ul4esSCN4kAui6
13bdvrmYXomA0zrhayzRelsoiIUJuKsktLgQUO2eGQeReZgR97IOJLJ71c9vN3OAjwK4QYJ6FglL
SbTc6J4o5FwR/wqjgyfZ6vW56rVVwbb+GxtDamRP4FXcZPBwChGMgWRryJ1go+BZmlh+UHzA5Ata
B25tHt5eWdEel3hJ2xheQAgsOoPwj9TOYmW8zPvoWkbwidL9K1gkytq9+XtJE51e054U9YPcLLk0
XPy70r+GLSBnF1xhdQCSUc4+cffqhHpY66T+tgKEopI9gCPynSqPSaNd4FNx44Knek36NAYELYJA
tysFFLt6BvfRUxYly4mQ9m0Vi/dG/bkXlfVlMPAD8pg4q+UOpeV/dz/6GotDI/1bnJzZp0gOZWvZ
PsX9Zyd8uegUUL8G7IboY0nLrFVixfYASbRlD+F1sWl07vlo5HklwpP4MGHbczMlhfdoannDbtco
F8xwaL8VnI0IHMw/dYQ4duCctIP4YcDwFHGrQex1YmaOnBKxVnmI2rbHJxRu2zFeTAvwS1MYaf7V
9RKGIa3iDWY5hvrCtOvzs53lFComs+Sty0tB92yJxxjcdYsGHVc19Cv/buA1PbEaI6HrgsOwLxDb
Qs7ZG8BwGGGxTAGMGqUvK4lySnO0j5IjHq+yBTrsSVVaMr70pLNSDIptsXwLNyzPYp7F1QKkZD8k
WMksr+iHRmrUTJPRinxC+f8bheL0pm4MlBz8LQ156DsfEHHLbr+ib0KKs0t/YPXWMMCabAT0tsQW
ZwE6j75L/tieyV4XvScO33cpxMafIpQmLmtxMQF/IPp3eG/95fJuJDeMb4OarBQZ77h/C1ey43N7
B+5u1NIKAYIxMzVbeXIY1jyotTdu9Rh4xqfrLMeCy11SON5+h4DxzjPmRRbACl5V73Y+kaNJJgWv
g5qRtF896co8t6bSs1qEU8e44zGMspOp6uY8CXnvA3Q5lHJbq8nwJOml5IqHa6u7I6KV/kSRW1PQ
iM8MltaKv1P7bh04+7b4XCgJpgup5TtH8rh+FAp+h7RzaOeZ8poVQpY4GbjQl7ebiCATtUxbqaYU
/gVYLIUST/L5rUSEPE44TsuIilYjxwOcj8wFCKMmunoTdAjHH9VJxzBjKuZep9Ue3cU2A537OMNb
tJ7uCvb59rleRIsA6o+X0jJ+Bj3np0XU+c2rdavheK5DMcnNLfjfczKmTZJV6YzIjC/0V0OEAgTM
BowW26PVO0+AtrhyIiZzLzXZffP+Q4a0iQDfniL0rEVz0YIDHsYA5keX1e95OvbbBGtdltd+CQG9
YD8fYAUl2MkaF/fngl2KCPkK9sp8E2/LNJNglwyDp4+DH2/NsPedc7uuVG6YSWOqSKQTZ7XVQDcf
15kbct3eYRFYiEbxYNAVoDL8N4gNJMhVPaLRls3ZTewq10UsZtPPFoUVhxEUMTy36wXJpkXlQuzG
qr3wxDND5lwzBtQQ62hWO6udQcBYJqx4PcTD/yAjcjjkcpbYQMixe0USA/TYu8SnLaoX0ajNdjox
FEd4gr9ioAJU9BGkqJEQsDx2aq27a3P+r+9f4bDN8OSTfwftLOIVCyHbPsWUDp2xnPx2+1fSe5Xl
GhoU//zfezRcVXUZBa42M9yQiHd5vajyfnn9F3R9Lv01PxaNkMPCj8z9zQtzUxd7/QCpjLCiWKM1
iXpewk+M2dPOS1fpnO/8xNsxJ+qW9/FZaU11ELb2FxQPI6qiGNi64OQQuuqbPmMZH+flXjwMEVTP
H3yrCGEdn1COU2mCK8Se4Virb6CWgRYSbnJyzoPQPSSVvuXzIIA5sPIfwDk+IsZsUJngdybPFNYH
ASj8MwKo8WTQn1D3982ZvY0cptW1kKOsCOAtA0C3nLj/1f84pw+L30BxRRrhVc84bOKI+a4hvYdh
k1iVPe6oFZi5LrWvHIyQADcWQj0NHnSiJDFaQFVkLCw+l73nw9n0sh3FWYzFDl7dzlDAJdizSJBa
ss20kPQpDuQ0EZC6ghF9lQ+MKY1rx39nAxNdvrFefPAqiUdTKCETkqf2GanM3m6hs1D5V4rled3m
2ntItoDq7FNyo0tOjUYF+zcW4BF//VBqxxefXJEB3o0NJrNmIDAKtLADC52nI6Q7mi3UpYP7I8ft
2MiBoA28UqiuCjE0SDzNNqYy71sIm73FBNlhb6ucVpvxHNRgeW/qgshY+UzeoIqEEPdkPf6OngL0
onp8f+Axs5ukIcvGT3RogAVbBLMeP8nDLWQFJGMHQnRQB7VzmXB1LOl42MWVvpqwfw1uWqAqK/7S
7RkKh3t9wywwrfVdaWPe7RKjIbCmACrpFRjCSRWE4LuKK1uuWf4IH3fNQc4H7GkZ4M7QxfKvs8Qy
ttJ5StpTQQ+1tG7tM5mKkpqIhtEL/m1Cr2IAP9UdbOMb4/F6T1ZJXLrqYPX5q+V0LqIv2i+2/TOO
pZ1fqW2TNllUZYAse2JU3fcGGQvfDZ8rfPZvFz7ye1cVoeDgbbEAWr5niS34b0f7anpb1fucfzqe
zOtk8ceg43x4j+hZY1RI8y6rAviQ/FVUDwyX4pr9HW8e/HlmZECJSxZ6cGhamDN+65yKE2mPrRXp
t4Bi9x54lqCwOrkhy7OCO8p93D6j6FdqdEX2GxeVq7EDNwXOf2JzWY2qYM6gfJJtPJ40xvwJMhOP
zfqdbFHeH1wHXUp0zt9+0jFsAvK5+10sjNvYIt5V9r/bC/M670hli1B19B7glRlLzXE1l0xB+uPN
XmdR4L0nO1KHE26/ivSlc8UEVxSCRrSJBwGTBPy63giL9XapOcvmO6cypzdAWCq+OtN+8jRdaD/J
iecz3X2+X79Q7F+2Xbdm7/2vdbmXXzJj19MjzqU0+4fugZcQ9tcTPMV8zWTkPDMd7P6OupojiX34
tQfZ+NpRqG6qNu07rTSXgp3dfWa60CL6zc3cBbzY79/7kQNxObfKDg0QqdVUVnDPDk8hnc11FMQI
F7r4OM+rlOwVu+hV3tmGZYDKTcqV54ekmzonQ1cHu2uIEe/aJBI9qTt2EenuNiuYZk2wp5RVzSnW
TWyqR7Ww2jb4Xai3QjI7QnQJcSAne1t25ouYt2xaxoJ6D2ovAWqc44U6uuD9MtOysMCyPAQ9LNef
s3h9aX5Ugml/zxxxHQ25PERkFWvL8jkXmWCtLh7WZ9xtwKTOuzW5WEZjfwCuQB2IF7yJghhzdccA
Qv2zaLZHtqds9UPQBQVXyenhVdoBRSbMGUbkHmg+mXmdY+3AWY4MgCqiE3aSIOy1RZFryh8+hV5z
6ngd/F9EikOl60zvIrKe24dNxe1lMyGte8MlLjyZA0JGi12CXkZ0n9hwi+2Q3nVyVYvUnFT+MI/q
y7RnQ8rXjYnGkdwXbMlQBa+7l6G4IPMStZcRmFHxA1/nZcBdD0/tQCK1U0PyLx2JaJWGPFJCDiox
HhKTQBMKl3vlOK8HKLfIx+v0R9eIlWnoEFLwX3EFCFTkINxBGG7OCZT6CxAYePqg+vubdCuVhQoq
2Nn3MmtAu3E934AK/cYrjULpmjBwgP5UAAa4Uq7Inf3veYvwpJ+QTG5OdeoY7Y5fCi8ii0TiTbLW
/vSK0V0TV9/IPk+2hG1GJVARwKLywoHwXI5vALnSprUtp+WOL2qu4XX8rBhoANrRiLFUxIHu98bf
AmcDX0HCuvO43ANa5KMuYMuvsxQ7tzc46+9Mmf6O51jxu689GqUORvjq6Qjm7qXDS8XgyXH4rtaw
EMBMcbPLSyxuS2UyqNSJXdEm/HE88ZAGiIruZ+YD5IPkhJYNNiAggNjfWjdfYnWNNrBG7hXO9VhJ
OZ2jyzlCwm18xl39Ui3kmjfqq11OSBxXRPyvtpjfTp7LmiaeFRjlRvdgTyB85/Nyqv0rUH4KKl7X
+p6nMd9qlKFTq4p85kyuJDd7P+lJSn5wjWNNGPZf8COkMgWU8Poiar3q9rHWI3KYA1nHE/ZDb++p
ZvVU8rmi0vVEm3bjFAd3mlBKeRSjVHNudz8KknNlM8WDHZwE6HuYwrZGXgoFCTb5SHc0awGSHeoL
mKkQBNi11jsQW5BjC+5v3ui3y0yU6vxZmqqGPO/F25tqz6ZjXCq4g/FCzsisqQOwqdVYwbNbQ/5A
gVNEBIo+isL4mMK17gaCSUy7pYitZjL1WxxIhKdVJWW19EP7IEtn0KwzYvPavux68gKWZ3KGEMkT
NC9uNCR70PU7U/hMI8JIi4Mt578uarxmYwiNiEX0y+pqF2c6W7wNUETV7+as49/UXY/8lTiwVUsj
T+SJ0FftsctZ9Va/jqPXZVlAp9aKekwkynBsKfOBLoDBtJ+3+BXk4JkwFdvCHxfauGb/ewzstqp0
xrJkyXxFhDUZ3RVEHDsI55UTKATJmQ5wKDLjTb+HDKspLT5U45DZvs+u8R1CaL9GW+Gqph+P38uw
paTHqAQUKRxphqhJyZPjpkrMnTKBr8vBkyMFHxxDlKRCpydgYkUFBXeP57PmwyPQA1GwCdYYZydh
fdRovw5wlPC5SOlk5jrHqhIARXF4euxoVBv7Aj4cF+EmhY463ThYogvag041mL2Up8RVABRt6rMO
91S8TJa7wjXxxcDClzOJVWSGKLzkdUYOBmgjyGYHQxCstVna9m/jXGtlvt6zfPfC4cwwDacopNYG
1fyloxVVYw/D41UWj7WAd5auYZKRzbslm9fUuZklhDn68nOfSn7THBXFmhR+9H2xyRIsFcVHO04+
d/23ld2f4N0BGGwnB3GXzMdK22usv/59uGzEkNoO7yc3yXtVrhruFwKCgiTg9sZpz2mZF8oZv0/1
JJaB5JR2/tI5hj4RyKGi77+mzfzgPbVeF14K8ImRp4ZejLLXIDx6ROOGqy0rAjLowCHDqo7EFzWH
1zhTfxiYh00thV+2MHIU/hzHC8zC366pBiPkVEZKG1IDmt64/qPM/P7KJ3N2OfHjt0MjRP3MHkgS
b3YDwcnpOiXP5+UX/iIeoPrtwZSsSBgLyxIEEXozbD5xzPMn2OJ+bVz7kdF+NJltmjHYLAj4RmpM
XpmEN+D1Orq4nEqh++qZirpumNTzEsH4T4RyOtohCOSKAZdr9mzNXCanlAX39OcMObvlQ3U5Cvlx
XR9WZ7KTrotY/xvj30ezsCU5hickVXjWqsIofKPRtPyfsT9hN1BA1SYG8EvQb5ttHl9wP75iDj+m
l2vZ83jJ0eCXAttkl+l6wU5o4uI6Q90Pqof90TUHcLZBo+lGxphHDb9fVp0MzuNxJS87ZlEitzc+
IIXbS2lpe4MZpMK9vIxaCumPp4anohGyKwJrf+JEv5n/K8/xDu9dJTgM9e5LlOjbwQpgXcijBRpm
t2g17XN2U+m92nAQUCNAdPNeEGP0SYCqphYjJI93FhZJSM6DZrpjrKuOddQIWAv940JEQ7ztHlJ1
sq4ZvnC8RVBSVx1pm3idd3Zgktj/raottoRcShIWggr2SVQnyTrgEliyNAO8OUqHzoayjB/m/wuB
vGKaBs6q+QT0FVJfcPGRVhjy4gkrjctoPtpHuYDFSuCXWaAI5p406OXVcslJQBGjL3kDNFWfznop
+OD/w0nC9mSU0xl3EaJv2U8L2FoNRQS3H0xwnKD4hW2lhUkdaA3SGO0NieQyBDkriLAHoHxOqjW0
kcsGpSWWg9ts94ILVoW7PgVS6TlraJ8hukc5Nzi9R2y6qvHM8QMwQrod7AcHyk2vEnFUiFU2Eh6W
lwjewKYZrFiuqmVPvyXg5yCOWVSsheDtI5VNEUQrdciabX7BMZ3YsJeqci/eFO8li5sqA65ogPa5
7+wxpq8iGzwIDGV+be7n8B5uK1I3h1OWH9Fd0FlbJX5kAtYqhTuG797FvBtcSa0F5XzTCnUcdRRM
q9W0QHyBjgaqaK8cx49huT0QMZNTs7qME0If96ibp405FentOrwd2/m2xcf9XzcluZeDTTkhJyIa
k31Cgva2HnLJNE9TMe4OE+0TTkhOXkMvolRmsLOusTRdJDgecOz9wDLmu0+5L7SID2cqUs0F6eKn
vyatqPtAPmJ76dr1NBky+XtjdqsUnITAUPiS8B1gjMkxgyNGlLkY4wcHZ8t9yC+DFOf0SfSv4sDv
ELYYiecX8EKpAqLgmx466K6QIN+9R2u8JzCSyawPoKI3FihT/XBZo+Uq1rtX3X2US4vbrET3ziRB
UXrQcYozGZ9dycPGknU4NXov5zraKkcmydIAsDsqgiIaE03xcwfs+ZmtR8jKUFqvZam9K6rR8Tuo
D9G7qX2+POX0+lBCxd8IlN8/ZVqeGGvmLL8TRkMwfkNLSqKOOmSdQ24ZeNBuafOMV3U2uYVZ6t8U
I1Q/K5bPxTBl4YnQKf9rbnV77MnxqrpKNy0bA5ag7tIiVSVpcmvds/K9xq76aVNHd7uqbcRMiP4p
OLB0y/oNc7Xsgm7HPID45sIvvMKgqmsoQWHPMAWHv4mnDhy4T1AVD8Tb/YwN/1xeubZVIoMkEFOT
tU/6JlEPLU8TSNbBiJbgZq+GY+xpu8V0iWRcDtuhZ21++BsNvqWdsEdf9fYrlegft+y1WXJ9jPc1
ozQ0gpDuyUeWp1X58dWJxioaFou4m6Y9YVPdOIBDdP2AJbuR31AJX2tZ/8C3V/RkOqNhpevjoxRx
jVkUyXPVLR2e0dGuNkw4m6zj3YYamW9qHDSAtiWs3BJuxRgmltRMhIOdzwKRXg2aY7T33p14Fqud
zI7ohThre4A13P/dh9rwTRdZKy6R/iizEcaQt4fxHgzEw99EUDViU9MhZMUiDBo1HhPCecvdxspM
A3FY+WBAAuXKub0ZGt1TA81alOqfHEyxf0uqGbb0lHvTO9QVOuyyDpcDRYspE7858dBoZ6X1ZOLX
Ue0zcyYHurCe0aUYaB5GnJH+SJK8IZpIsPps9sf6IPPXy5EQ+e9xGa3FdbVj9NqNrdo22AvIymyx
fA3vl4XD4w65vqbmWuNscG0Jih3ftkH9wgudYglmDK/6CVz0H+XRodk5NL1IKbuYqLQToufs0UA1
SPX+GoM4p/pp4ffaI+jYfTmomJhhFzwS99b8ziGar5OocLy8J9M/08Fd91e6KfA8pO1qsxNa7nxq
dtmwb01PcyQs7LllIySt68FmIObr4BHqgr8I5FsMNSe2BuG0qd9SYXu7ayDzXQyTV9h0S4a2XwBE
TuKuhIW8krqPgKOkPn6z3VtTJ1kvHPu0ugZ1kPz6f8IJe/kqlSVnH0FOABuCyWFwukCUBQ7Z8rS/
ykOS3J4uGA955ygAOoXmYUmMlU2dlBgM6u8tBne62i5kxV1x9R7+YtK99lI5YAN+2bTUwpQ1qM5i
9mtpG10a8FBofoTgPkqcAp3foBrobVxMA7j19/o+Ei8wVsphhtiLE5ZlNfKeRDZh4lsdwq2BeGsd
qYsv+6PY/Vj2M5RraujB5KJMXwzWBhded18ksYVLaqGwM9UCpsxshemFcdKpn5nL/0km8WPUbV6c
ccLD8/Czz9Lh0OGvxJW6v6S9QVGb21mzo9gnR+aoHkVjbsZS6OHs36YB6RGUz+ShnSPslH69hHf2
tVyUwVlX7VKc6lQdR7G89WVq4kUC5jh17aSJviDkUkWRUFPNwGRG+M7CPECjbM9CnLv+I3PZoVme
efQ1/+3YMpY2gyPJ1IDxFy2T1fSRwxw3fHWABe7YOlsviKoZpiC0Z2y101/ufsQ+ZiTHTJsYc1IF
xpqrlfaQF1x9bFWVSPMZsvbT/nHfzoeFDoU2JnVveL2GdmnDBXqXez+0IuhNMpNp1vyK4DSyZI4j
TkuRvcjJ77vaDipKWsh2fm64nfFRqkq1ovFv4X8GfP6wK0qWc8wqgusDEhPOM2KeosUoQ2qL+NOd
d6QR8tOCjSlEChQpQ3eyPqaVzIspIvg4MUk7rAIyYtu+6wY/ulHWXVt3Dhf0pyl/+ef1nYsbFnqF
G8xbAwg7yMEGPt3vspPt12XLPB22G7nOguk/S083DD1Dqx5BVibJ47wteMkwuyWgDx+tzzSNGcip
dtc+pUnnCXZze6j8lYW856ETeH7aamRcc+m7zHVtuD87igKwkdUkvL3DkDGY3P2Z8EcRk+9RUnjy
OPGFpTsNhUxidRA64MOp3LtAGWdflK7JN3E+qVL1q/u0UYPEDIaVLlT31/A40+0JgxHkFYCpUrAQ
W5VM0fMiM4ImfapWKmKoez9MSymDxZIXtegb+9+okGG+fwgFJWE0X7IdIPGl7h/jhXT/t5iQPDRi
tL0E84PJ+V1da/igKOUEDRLTuJ4YaTMUnQjOJ7B83HSY4a4+vNnSZuwcVS6qwAwICgb+1AZlOk+A
ROxj/28Pht2TanaSIrrd4Y/3ffVdMxCUmhlypgLrIvoIWkcRJI+SgTAf4FattjFmWKjshLnUb6i0
Mqlst6kMX07TnckvwlWYLo/eX5CXHNGtcdyHRlXLLpVRvSkr7dJM1eaWDGpzSMbQqk+XoFuE0/ka
Fc0xNTIehNkZq7xWwJqfV3OH9eY1cogo+Iuwquhaa66dWWfzfU43nNjDJqnpUGGaN4mr0qSTjelN
Bg3H2nk9zl06wYKXjrpJpfCiUKlXIMIVLfqCQAkvGOlSRgtsPh1sOY67xR40OeKsQ3OKoHj69YR4
5GBamdNCNLO20DekJjdfqxgYGBUb4m6P59fbPI6WDeQnM5G+AoxRdeBjU2kyuvitxMSMbDW347C+
HZkag6FfHRj4IjHOdNvE67sf7Y3Yas9aygXp6Jf5NO2Y0aS5hhuCTe2rDGSKSJA0b2qg42DpHkUD
oV0cwO27Cf4EkKRt7069i4s8KPGzlHFhKh9b3ZVeiK9UxDV6Cc6ww5oWLSuTbwuGlBNE96MiMPcj
QL/ce8QGSJ/7BM7yGAYEEo/inJMg5ndt6IpyLO2CK4qmkPszzXxIS9gBZ0UPmzgjC/+sex0trrwQ
6cvTXl05OJOxHi981mE1Vx+8h0iXrDI0VLfwC3oduLPyMXm3XXJcAZk2hgmjyc+R/MJPX+tjxxM6
uJcZcO5MThwRWuo55k3z1gZNcZnlWn4xDF41+C2E8cyMOUmf6gxa1Y00EUoxx01oQKeSk4kzTOT+
kj/sHhT4bQqzBAztf8JTYkIoneGzJhJp5EahJWygInOj/hml++qcA7ZMZ7ucw81YQBUJVfzakR5U
a2hkXw8QRQAmswGxv2uYaoGU0oTJ8F5jllS3AB8egeQLPHg4hZ5EtZrsfDaCQaptoxELhS75MbVw
3u9y9wv+HeIUVgyNvkaspHBAe+6WVGIgh0qz2T5j0fMcHAWU8WUvucFMMU4OYaOpdsBPme0CvqRq
QP6cX+SNJlJUnd871Vvd6P35aU+7WB7doAl05ovHnnqn66alXPENjN6qOWfWBCHvRSeJ0zVFykOG
bct3WKYUzJTMgv94ZiJYSHU02d6zV6yxxytBf+HwqD/ItKSfBn65AIEqgVgsjFHec519coHjpVyb
CGgMJk1KkVscbAmvcIQBPEOb/Cgc4/DKG2/3v4yDs7YxCiurG4oCHRto31fGU93GIbu5rd8TDplQ
kydekA2H66xFeuvYF9fHR45jO0iDtqw2tveJwkRJQ+6yqYcWlLiVu/qP92j2zYP4yoWNKJ73BGTh
gXjMsGismVhxNnnKK6G4fRQ4SbiguSCMcUpwnt5sHTHCN+xIivmXfCZDXpQlF5fLcV2TDqaltqdm
KxFKRkENMo0uurtSCuPwd3OgJtlp3y2HTMm5vZV2jb2gDxIhBDaf4KjWEKCeFzxxtDGGqIbNjubI
ZyLMzEsPESoreMSbgVPHdQoSszqNmT2d7CTOHYZ7AAOwm7nuEESxILP9aGIUDkoGzupOhegW7cQz
MNyqToCuwar+JPeG+1DsEEZNxAcu3SMNi0/9iE2i0yahpInSR0P1VvW9G9KUqFM34MGCRfNMchn8
O2GWdZVQ+5jNn2CBvs2EdjOCyvDbhAWxYbe1YTBK1qQ548FNrQLt70qw4xIO8IuGp5PYDQSGeE5n
t6eKl0br4ruFnIiSqGI9YpHbq1+GZ9LjtIPz4N/vw00IuIDI9db3d+6CvzORfzFFngkWm37Cba55
9V10jr/0KQfNAIcPmt3IGOY5CBoRDtYhYxQYAYDhwBRkYh82SWIGiX13wrKMBF3cMKf2CCDkGCT/
gxXAMd2IY5NH1n/cLzJJ6s+n/5+qXQRBuGJ56EV1IOy/Iq/C4bBPew9N4BdZiXFbsgsWPlGwUryQ
tR7vd5BiDJyXhprRh0ke9xEze2FC4PnmQUZgZI5IWwLE0RZSaH/C1dt9T4yVKIBv3qJA4dkrGzwW
lJYBnbPJV1tgyrtYzEG2lmtbBZd7sQLHgDuMdKz+V7e+DZrj6I3Qgu4ewdrLXGQLAJ00A0qRpm9q
F51sikx32RjggVHgP4qpYhoFxPYW7gtCaWJqEnTAa91eE4jjoISRF22zDGdgw+1k1CZ8SElv+xX8
tCJuU+zaYJu/JsNhV3Nvy7PzR601F7a04+tdhIVpvGilmNLefOLvTTzlvFlFEUbfduMpWQVNM1L0
BqyNfLsCSOmA0DDNnFE4vlYtQ3GNRy0tql/wmp6rsFIcRr/NdeHOfUylsErzidQf5s+tcsNNF60o
wmaXjIK7Y39Gj7K4c4dVVg5tB75oQIZvaURtV3o05abOZeFK+wiOCStz72OJtXDFl47dTLAyZCXr
SEzw0bvEJ4a63gV//T9Kr6Un6Njslnt296ArDYn35X7GHDH4ModDXQJy0x4RGTUCpDKQbBRjf9hv
4gdi65ZdhtF/Aw7kidKD8c8tS4MiNic3zWJ+za2p4O+RCnYOZsCUdQQAXEUA4MzeZgsBndOnjU30
ltlUJPKU7TZQkKDmwP4PJJAyXg5vo46QH/cPZ0/SdG47UMVXku49MFuG9N9X6Vao8sIJcIOgMcDf
secANIcdATlGAGaDGskHLqiGlJNhnJfLPMaDAJsSoNEcL3WuHGCvOj+Lyjpp1Fiqnl5DSIDdh3o7
sWqLg1g1a214hbMIFLdjzgdX0hA7wJZUyCwr5cBUYUx4YKTadL2RbQUTy7AgoCYzJCd0hXo3nsVr
ha4fqsElVqBsOVMMj45fe1ReKo0ukRrbhdDO3HgdO/KDTj/nW6WIJG2eDuVPELn0Aq7tq3q9Irw9
+GRP6rgdETa7AryZvCdvECXsyFWJ6kY3jrNYgbP5TCRwCca4nPDokhzo7+OYO7XsQ3DOd6G7ZVVM
NdGtBHn1OmjHEjNyqMNaDoYfOMtyclzISpqMAbffHvMGBqfxU9Lqlgbxtyt1Kcy6lySMiNaS+LeD
dMSG1Pd0bGdo70SjlDeEOQ9Knceu8booDbaXGs3ZkXDN8W7GTjcGCJcJOK1jdH6J3kgq+FBQAvCU
54G0pF1UhiJAO3UgxW+ouTw8X4p2KK6zzhwQrBNLKgbaiQupaY6CSEIRbP9eBXR7j+sbf3oRAkHK
ExeDu/Uxh21qT+n6BZapTcVTfyRsNV17Tl2oi3jMrm2F8iOVssnLhZ5bmgDIuOhO3CLnWQC1JYDh
30K0ZI9drQOgRtRp6QFqjaTkzFqm4bscXQ8i2YeupHCFgEAxa7f4S0AverkBlTDqngZewl0RwuZk
owE+1cSDqerchtiszCNLQoELn3GQKpB0DF1BVtRJZTnpPylohYZPDllwaKuskcmeKLodrrp/gan5
sKhz+rfqcJ9EzNZIgz+4ZAaQE/RGmTBlXyHjHk2dS71lHyo/r/HTJUOSAjFV9xDYR+eahZ0TNjpV
DHl0eCzkGJ/1rfpiz+qUErFnZGSDqo6RzRMs9sbz5Y5wNhuX+h8fWo0Ol4TwnvpF7S35z+VKjH1l
6bwfFIx6YBBUp6xJfyM4kPAKzu1L1dlddqNxLbIlQgIdrmr6HCLjRvYQHPOivBjBXN2ju9/6YNdn
E/IcJXJzLPyurO9GWBk9mrvv/m9e/QYtpUMUzG4jVx2bS13T+gx6vAW++JqiOhKSVn+9rY1CrWZ6
ud+ro2OTJ/eA+kgAYZWuHCFBwUaBuILYb8+Mql0U8jSxw4htF5AmvhjvpI3TSeO6bIF/fAeS81Zh
CQBxpeG/SXmDEZxxVQfRyorPdmjbcyMsIw8VIatDTgs4PVUAwI293+LT9s2lW9eWmzGmvu8DEKAE
jONmai/yTx1QMKs2Z5dkqFUPx1oiI4Z20ec+0KGy+rAkSiNdv6ikaYlNBR+wK+W5h0O/Opf7Gtz4
HQstU6hvkA69ld/1y/beyg0wrpmP4R03dV+dQhQZx8Qz1evxlpyoLk+ng/5Cc5Ihf6UrdJDqPmX+
jvy210LixHyWvaBhJRVSODOQjTEUEfJZv/8MxZaPaOdaZfqNxC+5ofvqIBlFWt7AOg/r+kxMHBox
KpOppLlZdg1lMqHjSqeZZCiU0Afj6sTp9d6NjBQRA/FiBO/bbMQuD9CJocejz8OA7y3iHepzvr60
bVgWMsrQ8J6W2fb9Hb9RtdVZIW6zPOPspOgjsd0HjRJHZ25/GuBU8HkxX98Cak9sBoZKoUs1lXa6
3MjwdBNsPwwzb8Dag2Pgk4wCjUNTun6oy8TPixYnAGQZsXiu0mAcBLInnsToNCNBwSaXimu0zdZC
XmuJetd7gj6bwyJ7sCcDDNFKkFupL1+Sh2w9DAP/QJLdnnvdgnYM6iEg0FitFXrGBE4HCcK8aT+m
DxXmlUsV2B8Ka/QJpdFGHAKRuvzOxlf8rJqU1L97Znpe80YDKA5QkR3HOl+BDbyqJlMo9BtqM4TQ
qPzfMvNqJLr7AFVqffGbKkKr0TQYcoPHrBgYjixLzAozdPkNXcPLQCS41JzmL622wMqXBLG6JL9z
X2zrpkK+DTqB/febqLTMq5HF5bVDJlC7UassHBmRUXQAUtvRMEujH50XTCeDBOrqps0wkirC52XC
guxv7GZ8ZAWh+aGbqIBmNdDrmg7ZcaPbFEecppSivdZGuF6z43lFpBpZykpzNQPR9Yeezi/BZPRJ
QYj6GvYa25ZjJFi+v06NrPR5qj0hEf1wAucNcQnSPaDSFPP45KxNv7CkDrjduIjFaCqn3hM5VZgN
Z3WhfTeVSSfDm3ZvVNwTU7ZX2oM5cqsXC+zGD0gbBgzLpL4OwywxVlNRVUSGYGPq3Z5AX7RKfsfH
Ka3pA8Zu831PSnSCTMdt44oH5qP2sa1yVOjkFoYKGU+J68kn8aJoWPmzhEaiz0rjRNjZWNdi8/iB
+AcKPaAMiC2R7qHAwpxpNJj7LPBkMXchjNzeB0ZcdZ8b4FKXQ2MHjbBCkzOJTVbeB/GFPrWh+rZm
jKYtuRhn7B1+fKpcYXdPar5yC8QWap1xBRn2D8pe9Wjr322bvwEMFYdcBzxhFbo16k2G+WPun1SS
okErphCKN0xGf/ctGTiM/FjOm4lhd7n/s3W7/u+oQGDaKM/5M0TuZtyU4PglHVSgbZmWbp1zapx4
y32kdyUxhjjsrZr6eSXkkRCD2hFLBTSqfymhAja/GJPb224nufBXdRJKqiPpqgfUF0qdTf0kw7+z
Lmxbbs0mr66rhU/WHzq7RffPprypOV8oMxLgUB3S3JE9BrJrsaxqUDWX9Wz+EcCBtOl5q+n80RhV
5uR5pMMlDsuL77kLFy9ApjDtgKU1dU4HjoArfbRrv0jRepaWngYuRt7rBmst/rySsCw2hPZK+z05
2613JDd44gAjIC/CgWpRzA9Tk0NjugqUemwst2e1qAwJZ3xAkcApQLo0+O78mfatg3yt0bdK88LM
Qp7OvMBE3X1Sp9vuaBL7TATz7Qj/3INOjsbw6BL1w2kmrxVadHjJhha17YJSDGTey6JEApbSALaJ
cK0ToGiLHUzGdhtPGSzNCq/zCLAPfObqns+2s+dm7iFoue92Og2G//sCkOF+lv0xRicvQOKBVa1U
uUm4ZSRT9Rb9hKk6hl4XjME/h5VLz3OBPd+xyRLe9bFTy3Hk5Fth8QYFzs+d5MnYKkVvR4hr1lyN
iNW8OpUVZsnO0jZ8qs0mXYccvvEIheDNJ0moDCWYICDUVaqtSyALI/KGPmdL8Y0glQdlUyxHINpL
YBrE/injevEJHMIouizqgt2X04ourjtOAboOODp7QUr9VJAzKse3+y4XK5cOaruV3ZSe/DmGnZQ/
R/35t9JkTvvSBXapgsXXfxdeiqMTBgVRGHw/N8/0NyTeE69dokR80n2pEMeXe2d3lYddRAG1Hv57
gQ1J184IFw6gJfLxjp7VGMd//QavQufY1X4fK5t38SCei4nFlcdCIPDYPSeN3kNg2QqE0vFI5prH
5lQ80yyENm6VJ5B7nS7ldhsyjM6onWMVcwNemtr8QkOGp6Xh85CA5JHihlJja01TmvCbswUdhWZV
BzOTsFmdDFLrs9nv3NU72+X4tmb0c0pVMO+yq5hf4Y3kTVEdh9qfze1dMeFvqg2RiZHAVDcIawQj
iZWgKOWAAmf6Mqu+Joy4oUN0vmo/Cxtwwbrv3/WQVAAnTbAdWaA48Oyv9n3iXaPp4DA9lBVuusWc
njGN7cIxQvKTA+MhYo80ILPr6Zm64VAE/EqVvfU70ZzPD+SAQihAihdSIYMVXvtXkDeaU1kzCLtU
PidYvrHKo2YIXNEjg1nKNOOABVPBMruda3bZE/obGiRdjt64yEG2fAZWiDg7QFqpb8jFfCBZdJ0r
VhChgmhzMooCWHW1w86ixvgLoLBVZaH52ipzbCTRDKroV6GJTZ460HrCd2PuqbcT3lLBs4tQ6CFE
jgSB1whqeZY3QDSjrCap6xusoulRC0ut2yZQ75o0c/PwMEajYfrtBuFN97T1ZPul+B+FPDiSPy/z
B3x1jGrIp2YXmey7cUWb2EV+jlDYcMWbxhklyL8/EOa7vl4U3bKEQdNSzGj3mS8tlpScbk5x8oF7
1qtKJK8ECigaZ4prWj5HbixjA2d/ySpRuFN4+J1qareBBQj8SiUxJLMeYtkYnF/l7qr7x768a7Ao
V1DAdK3e1jyuU5atYxatYBbkQRO5KdlgnwPie1H6SeDBrso8NQkTk504qsTHCGi8/WybZdPyiwVa
ZpGC08nB0G5ZfUta5R0YR1/vdYSQUvYn2Vs9z2mWOoF2LSrl+8KI//UMU8eaVspH9/R1MmFeWzHn
GUkZOkCYVIyTAcJz0UoCYyT1LhjQ0u5sEetn/AFenO3U6RUn79Cd1ny8KTvzLj4zwY/iAub/fX1v
qmIMmG9p3XFKHQfxeGb4kJKfM4Yczkv7NsLYKT6W+lI6oAxeWHxRPQ2ZpQw95QQNixs1tKT2kDUr
HulDJA8Ls0IDV5mTW3So4JIXR7vG3EVYdcFpsuSFDLH8wz6Pg6po1wTWV6vki5x1VrRD68tlokqc
axMFI7WUPDh7Ln/z0Ig+s0wjPyisQ6X9v+jpXIGmcPGPZf2EoJjaBwWhJE+dDSTXMD4eXS8BWhUJ
6FNX1wOP8s6Nc0Xq0e4pa/qTZDJmpPGBst1x9ZVDQEWDJEBGYWIXvVTP2MTmnY/VpEbYo4p/RzZk
AOFC8po2aBpNh/3plP2AhsUw1fUsJBvWLuvlL67FerpcaMfqN6u7nD4uHUCxuYzxQJoMAEz/LXOc
RKixxGDDsoa5jsXCnXf9Jex1LAIaiF0IS03r100fQaUVkmLv9vCf37EhUHeiQBnSooGMQsAjYlZ9
MxHebsP24BXWJoLg+NrP+X3+7ulBpaRMelyDw18gJGMHe+8qFDehPmmkOFr66MqHqQDw0yaQda6d
1yXB9VNJOGhtp6WKR+3rti3Usp28jpRwo4tD2gxWTk7bi5hdpfbNZXmrw/bgK8hQntIj+ShyDSvF
N7l8x+PkxmRnzdaZimYvP/aDWwzNfpPv/HbWy/ix8D0/p+sJRbZ7MoegPvbffGpLk8eAknMsQXSH
8vhWyIF4oW9KiWNELkHDXUMRd37dJsZa+apJmJTcg04H/BigFon937hBV44GRKqUK5QU47W0EgJY
keA8qgDswuuFSzpL7b/GKkeowDpYTme7cVfmrXNofMScz5qyKV58pYsam8nKjrU3yfO6ORLLlKUz
Wb9zJ5ZRRh08l27zQbChDKHqVK+5BfaUhWbRmM29mAlW8VicIWpnEGfzAV+x7nfajr2yQgFgNxj/
P501pFjNVCvS95mQ3EbbfvN+7fttPZ42NTAsxlVyTdFYalbJfab4MfRcgBOXwjE0FdkjXhHbbEkF
0K9MtwE/4AYYo7BbDNg3NpO8jBhp5diIAl6C1GbCcM2KSNo8RzaMQAkTh3xTRVnMLGyYWndQLDdE
ufCQqmHeEJhFta96T3/L7VAHb/bhzk87pUJiRj7AR/ybVzJBy0NlgY1sWSjn4FDxKaYX4mCuJIdR
bIjvCSXkvo8eFI2bHnRo+QZHXa//8YgSmZAETNwfr95nU8rwnFYGJXpx9S60e4if3XgU17UFtfIE
b268/tkw6bNU4Q55fFMjN1rNLcZ+7X354aept2Dh7VYVUtyf9cFo7hNx5s78JsET4SqITJk+beaJ
T5cH4NoW9lTqcqDP1gMazf8x1YMhbBqcs+JfMFdaHDsCOemeX1aM0GIl9SgY5KSEotlzRWZcC5tC
ULfX7G0DJN6mOcIrFRamEvslZcvJ/Kx0wqRJagOcTe/6Q1W4CxatxQwCQoy+FOCuDGIhR9vtc+WB
+YXWJpCd4BnqMaCBslrOmmZz/X05Pf8XbBw6ZBwaF6cCVOdoS269J2iMeLBxnZkdi6z2v0zDSgLF
6vF8dEEwupvLsxRzgdv7PBsA8aaM8q1xkanKl84ufuKzovclUarPU7EhcnHcSOvB+bs38ql+fvbk
9MZsOExv+d2zfIzvwFDokykoZWeUTDgBH4PdTSAV6NzmKo157NbnIKDeLrhhqaqoME8fqJ+z+3Wd
jfLvtkor7PsTSxUSaSLY8eYIjVs1ymO0TVxiXJGK4PoRD2SnRNGIBeTwL4OeOyYJl2c97lSSgWmD
uO3praDMUVtVe0vmux7MloG1/xo5XvppZTvN6rgcSajhaAGt7fB8stFj32x+Wze/B3xIursKD0Qi
OkbEQC97xgtHpn1Bdw4e0N2848RHyKOMrFCFGV+JKp+rIawZlgMEAy0JwIids3F68qwNhgYpW9Xq
0oa5TOmOB3CIVIT9JRnymnYmBrgeFZw7fOT9hltZ5Y7aWrQ6j7Qgmr3YBV5v/abfrbjbTOXRH0jz
RkffOVKXPUbXLSCRG0igTnSTtq3+3srNo+8AzthaQ7v7SUUO7gbRZLhT1/5pj/sh4O4GPxYMCAmP
0TPNvc5z+0/6+AVxtCmWOgAjjIwGT+6A20yHsEJaynTzveX/8P93VOocdGvwa+6MFY6RDKxohdP1
c4THo3Oca2PHD2KgL/5M63mDfaAbokEi1PiD0jJUh0EtMNWgXPuD1DwYdY58ErNrnz0jeIfozhpO
c+EZpPGtFtFjlwXsc35G6FGlhRwxkzmaVTRupAoEw2TjTnrsJ+IHJ1y5+ZztE7C/3R70gFr/Wah2
2zNkIFPiFZoB+6q5JR03hn4fTUntBiXb2340cCZQ/3TPccJqJUmw1NsUC7kF35x4XLmquR0rbYj4
aW7hNr2FNXppiULeNyZQ6cBHkt+E6YYNx/Vlxr2Kewq2NM7/BQcWNTLMhGSGCNPn5DMGmWAUSK/7
pB9Uzi3z5wI8ifn+ehzCQor8HYk2iBQhwfOPsHFiFKAigOk+/6V/BKnCVbJe45zuoOmqFgTSiJx6
1gKN0gZl6uuKx7cCr9/FMwTUjRgSWeundrv5YeyJ+OiuD84t+3kO+aNnkPpgW9S+GPXvUOWwbhTf
UyqiJy7BHoSYeBb7RTRNi4XP8KhP6PFM15Qc/EiXp+v5qGcEYZb7yVvLPTVdGZVMaeI2UUS3Bc+L
C0AmeSr4/vqggUGfrC34nFuYRrAgFCJTvJUahXOFlXN7qtqHdDKSaOAerSvGniq+ZjBJoAazSLY1
clDhd3IZa3BL711+3j9YYDZu6Q0h5V5WYdClG/4kxLO9UI/Jr0RCIBwU//hjqloMoRAYSO+tLNkL
UmO+bzGlEhFgsjWElMhvuXo/EcxCZ3KVLetUvkfyjHkVGUkOXxxXIQd1S1G7uIqfe5x61cufA3oI
YD0LU4/fOtpeMoGq6+fmvvhR3LzosmCVTrOXwHxGjS7UOug66ZcSYiZ+30nbRUXAMFTY6tI/aKJ0
KkHyibRdcYLsNMwYu7VetgE2hUznMs4s4EjydjSKviBxNhR0zqvco3MpBMejAr0k0P/r9YE9zXHl
uLXtVVth2Dp8/jzDPU8m2uwhJmtWUWDMJDiqURWwhKvQh/5P20wUCOOv078WyNzHHCjCI5O8q3mq
nPz5Y20QC6H6fkNKg3Acacjt0z0vsmesepXJyaNNjHmURRugjj6gZoSCYIHTdZ9eQY6nS6bGJ/Nj
fxyUCzo9jS6ZjDBCR0Axu10Fl1XmLLL1tlyjRP8in5cpfWq6CvzV4Fa6QVt7PnGPqwiCibJ4qU1E
cQ1iz+oCm2BYsuq+LUBgU9qorD28GAj06meHHDLWg9CSXQex0TUJsCIUV/XrVpsZM6/1SghK6Gir
WM3mMkkc244koFpRkcPw7RyTdiDfRDrGWHKPpTgn3yrr+ZG+kdXf0l7pGUlbpfHRfgNkXNVa7n39
3emKuAsCO53RZMYb/rwdcQuZ3OFljbDdF7hb4XZs3914XthYeoWiTUntdO/cxdHyRvuBrkshuybV
SX7f4k9RWyuQZkgFLURk7vWjvNp4rPL7mY5xpqSqtWh+OBcEM3qbUq93Y1Uu6FMbKP6gj83/8sWb
q5aZ+sf3rs+oFz5So6gMraSF2Wb9maqfzNHRq3ZTNCaOoiJoj9bV/eqP2zu4c9suMMkLVXIjgPNQ
9A5YyKyOjlX1tzjyjWquXEX03+4d/fougt8wh0oDGqQeQi1rhVqiIrj/AmmuWbZHUV7ZpY7/7yLq
15n5XsKoAFk9juKrwNMHYbPs/Bb03ZYCb/XM5geSYbvNxUjFn27/o9pTn11E3K2JYv9AdwX6UjgU
fKrLnu2VqThDRjSQj8xULKyNM6+3egOW1ZyeKGbyuf6ddHDF9ygoXSZ91bu4MmlNFlmoDb/2j7dv
1Wv19XhDCyikRYpixzij8UQ5JnSdYAR6duInZVuK/cSxHH/Yki6gw6ZMySMVTzqy5mg4GQI7U432
Ow+PFi7khHSXFmdwB9si+GlKlnvYc1zWYqMV3tx836g5E3Wkt5Ywpm2JLL/OkagSadwDbF/snOaE
gXc29T7FkN/mh/L7VueWC/6vGvQ+Bqx5HSeJZqSeCrbdVqxhEZOJCKjqEzZIPPm0NZ73fXv4Lspb
xyCBywmEL94gLV6hsNofojw3dYTBr2mN0b/tnjujuSiu+UFqYwuJt2sSoa1E89xGbyfMuCzXAF5x
NCmWjQ+yRg6b6Hgw1qvdJ6CeSjRHd4PJPWvP78zejT/NuXEJ3DIq3/Hg4NcBK9WvLwy4x0OMotFZ
SktHGs/zUCs3axFeaubkZ+5xIzCVoIS9zBwqYxb1jFhwSKzrGPKxLu5GvKimrVBTkkf4Lube22UY
fgVBxbHzUMCiCR8GveBzCVh5luTNWC4bNmG54SXVhOaXCzVuPpFMg+6oiJ150l6i1zbH9RWb93ge
rQEGiURT1wA9iT/UdwZykr1kXK2VJLa+QHMSOUpqsvb3AYv5HGNP31wTjA2wi9YC7r2NC0Fk4vyr
H4Vd0v4qOywWO2wMrILg8c0ULWR9GThYkznsFEcwAD6IzkzMdEVEsQiuANtiRyxYUeQ1G8JH19GB
V21iU9dxC2b/y3vThdb0GEba2avNLqrazC8VIvJQG9yglqkCHT0EU3xqHNqM+0+euU/S4RQnRpNw
MrUdpj31eefyEBhqxt/olSLYcr87qyWnp0OfIOHwmDVnmBw6yPVpbtG5dAAxBL1F5PjDmg6DKaGH
RoNpdBrGRqx37BIM/skMslj18aLcQ2lTe+y6cMOkhd6xHKuBpHsQ+evF80Rv67Iefy8o1D/G/PkY
+ub3lJuML05Brgqj+j0nSvDDb+jsg4VJpVJ3305rirG872xE+OmJ+c+OV61BrSVdR7TnpkfRfylv
XUmveWJ6vDOInsToOJQO0KnjMm2+DNP2fAhPGgSD/BIOecr/lulhxrVx4i5fmt+cRFPZ/Xllzyaf
0U8XPylxNVpttKmtKpvGMivUsH8Vm0Z1D9W2rNeCT3BPEiEqrwzpQZ80lSSStn7nM1uaHkQxse3x
FVQQSxomerWlbAR7LdYdZWntxPgnhYN/LLr+xiiG613+FOlJnmvkUCAGupsLRqSW/tJSVAHAWH4O
j2mQ43jVGf9iZYVLFizLF6t6Xv9XdYP10RDuzyn1/PhyOEZS1NMUMISqj0ujvwohQSe/1vodau9Y
dxzpMxoQbIGmMIoxvPzeUyB/dZK4m9zM00RzwTQ1s1MCq6VWNWdCPRqb8IfriV+YGpTfEZXRlBmh
qFKWLLmlXbWp/nKRw6eIPoRCI+q4kVGln519Nxgr31+Mn/faCeC7OmZhJzMdlY2YRmGcG4mKNpwK
IupDH11gOBvG88fWzvd0GU5W/8UeFRawvefmED8PsNQZ0kOTy+61SRay+2P3DZ4PmeJ6GGsCigtc
lqk1qVaG8KZvTStuKpxWMafHLQQCbtlHXqhdSqTdUsdPvcJdfTeUEIcJIoiwMsrQM43hIWiBEmhb
38TpljRuEtLZEHSyMip7HtwWRwRPc+1E5T81omEiB4o1Tc0OrZGflKW7+v9RP4v9QG2brhBgp3mg
6PwgT6IheStmWVJeCXtVyM/h3MI0vPJDnjP5IBJcdm7Wu5pVCV6UDbQhkQfzsKcBLItIkyx5IuUP
AthvsT0KlqkBTjSusjGloid6FWCq7NzHV5JzmZuSWIKBj/N8LsWPYLpyv7bBG6IBIN4CN6JqTHb3
sImw7NCIcDRjsMIS3xwouMmnGu5JdoDrpq27/k6PEyGjBG7SZ4MJ+xqSgOLtm6IBJEPsO+tpvF0v
hYPrqz2RUXJDPMUYK5dmjzoQMeVLX6HxVKRBfS4Pn2VeMHQOA3ArFsJdmOZ5s5yTY+I8rvcvg475
uCvgs6+sOGv3xFq9zTgJmFLygEGk6hh7f5dJ5jonPNom1deDq904Yel4P2Z9ASkeRxyk2/xnx5zj
Lb9VRZnzTUF8VH2GNPU3by6okurVb79NghIFAQcFMxtYSOEb7MjyuYxcgnqCynJXNEiDlVf9+ecd
iyPwdHc5UJhHuDKMOSAh3ca3JqlJhD2/FrEmcKXygHHRr40IaGG4hwumFvmx5AeYR8Wl+f4V3oy6
oUQftSIitDQmmXbFbqHxh5j5wXCw/TVVj+8pX2tWgZ7grCVaHNDFXx9VTvxcD3Qvmw+8FoL8Qsaf
R/lzs/03ARe2q8V5saGJ/k9llb80hq6yQkiddrkxOWqzyCE5/AEW+0XU1Pr2vinofT3WEIZA1lhA
xiEx4HHfWonZGpMznokIOPTFlYLfoz0t3i+SO9ek8F82YHqkix33FhH5HmoREatlwdDHZvYQ4he0
YVDUj/udR4W00nEuKWyrgpe4l0JPDaKFLh+Ysrm0YW5dJnjNXPsaNnC/NtOwcKc49M3BfhhOFFCv
TFiKYLWqwA9q4wEFdYreYwv0Ik2OuiZjxpCLeFcUH7sinov5uZQJoMs8cuCKeSSNelSQXmurEy1X
Ttd9bHQwl/MG9jR4qVRqlzOQWTQ4zSSQ4DeqZCTMttWWDr3hVnGYtxQrFQtoDFojmLvOgAoFe4re
CGkBmhp70pyIJhZOWeYcKBUSPqzSY3vBvi2KrpbO+R9ENNPjEbAc4bl51sjsxV2DzXYnfIDpJicg
wIkYHypxFzcbvBu9pNLlkHuWt17FI7n+zwhXruHLrmAHID6LSv6pd5XYKJ+wEIQA+d7ZnwZzwFcr
4AgJgc6SL8qEZIgpgBjIbJbY4YV/0m9stuEI4Yrc6N7LUtZ5QMkKFQoBaWwVKFwFX9hu+J83tBzX
tbFIebvWfBE67G2U5XHW99Py9PmlV3rV49DmIIHuIAaRVNBMknE2e1h/9w+ydPNE+YO6KMYRBnKC
Gty44iPWNzNLTk6a4bESD7hpYUuaOVo7re1f+SH9OoOAvccdQTxIX/HnnQWAAo9WA8JHkCAUVJ/y
8nM2btDH/GOp3ucJovZUjiSieBMKriZatKJrpWtKyods2jFrZCJKqY+bMMiLAMwl+i1xl7QfQR9P
k9+TtHNL2M51wWCcePlXN173PHOQypxWwMAmKayi/O63OG7XVyO06Qyea6CL3XEO8zXCX+3vXpDz
lKVF8HGljI8yc7R7FKsfRsRKRVLo9JDxqI1mTTSji9UVezni3wFt53UIQXqfYN7a7aELf238rVyf
tlUOL1+4EtY1URjvpqQezUWiQkK3Lql85Pld07x1X5ZZ1I3aVfTai33V+GP58Wgeg5cLVWvpi3gP
i/EUSw4K1iDxc01URhcYQUw0vVGzpeQLFnY8+SKUa1JmY5kuRJdbN1oKVCyGiqDSKKQ2TaP5fB9e
dXF9dqUZ71X9h3H9xSsCBYUJ3XYY6zH7y5ntb7mgw+esMyFRLfNkdMWQdPuvQaavig8tqakFq7oQ
f8iHNIIib+9KNZmK4pdfI7ZJhXYnguzVVSXdf7grdeU4Wl5aE1cQNB55kDqfF8jLbzB6a88gar7G
Q9+KQvRumzNzrDed8kGU6E1qZileyrKyJFTUkLkwR12O16OtPaKtCg3f/uw1wNC9oTNKfDqeYCwR
4nit6THthPoCR75ObT41pDYE9o3tCynB00gWae8iMK/3IjtIqJUsx81d0vExVKgvdmgsfDjTSXAV
hNPmETEMHfNW8wLeWInISJ9gxVmzcL6sfUUItePmc/J2Q4xK37o2vu2Q+WGcprR+ropO+vb/dDnI
rrPy77vTB9UjWcEBoMD9tlszikjrL1LFIKH1E1CFURfdTSz8CEaNDIP8kT+n5P75teXKmYAkF4+V
oD0Rq4iDIwZt/18AFIUIuOowy4BN9hJy2AUTsavsgilvXzuIFt98y98pM/7kLUE8mM9jy0oGexzi
lS8v1Sdyi9LgNTbJWasC/ZkNBSJnwVYjU7EEGcWpE57b7rd2yyEwJImCv1dTe3wuOXvcN5WOJrt1
YnFnLgiK5jeJ/Y6yaNJLkPzd2zKWb+tOmZcN8s0pBXM2Lyztmc3jAZ6dFAz/KP3WZdvcwUrStGsn
OXTQZP9J5Gt/vfOhLfV9DQw1KT17bq96HbDb89iNaAIY7coxhGC66nra1lY5lfSoYH4h95SfeKQ0
VdbBVm+mcrfLcLRNkjS6vLCiq+ny5MZZt+I4URk/kyRqGPYWDNGsWYdrRfiHdmntLBv/o03nIZTp
2tB1zulG8rjt/YHuhHddTZ0feN86rXCiNPSguJ9QjiHsKtWise9ePduSRXOjeC3BTZ96tUvzJHUQ
l4nR63oqQcFAgIVhmc4kqBfx3vTytBtTb5/mLDTwCx/OskhlHd9qTLdwXrLaZkgVznvexsY/1Ajp
TdrBPSFDyv4MD0+A0TeYoIDSGWn3tqpBNn3T24lXQAyfPrYfiIao98uc4SWW2IgMANER5j5B1g9X
YEkeRaMo8OWyPRBN8qa2xxCNUqPuFhCwTE8Ghcuv+K2H1bjR0IDz0+9QkNW1tRNEp2Om07IzSWfu
lU2DafznrGXrfPH3chhDl1gFW+UPGJPEWC18UFQm0QFgherl7B1/I6qMQfAGKemlVjhpUP/pkE8C
4uzBRMSsiZHbgakycyLMndRHGXeeK0PZZP/CCXX9O4t3PwVZqI80xsaymeKdt19425dZ9BOTmzT7
OSo4HJXUDaPhRcczhSUTQ6kL7lMz3zW75ycm3zA3iMOOziyR46wrxYmpPs3OXCO0BBpjwlj/GwV2
KCoWKlyT6OoeugWujrCDoWGTych1qofoN0GgKq7u8O72p7Xe7p90bCCygz5GIPrMEHFSjKNyBaJV
cqQua5nwwjasOsZ9HqqVsg5sr5ogad6D6AtfpbfD1d1bIFnQRyApB/tQM8FC2C/jLrxRvvI+MlZn
YtfO6MPYKyd+R6gUlM/5EDNzpkLSviilRDLq6oR5JzOle5BvW36w/eG9y3Ph6rAXgY4zBOdN/bYB
YJdOYvPeDbW7JwmWAuyW9/jyuO5dqKPog/RxR5Q8xhelBxNXapjZGO2BkFMJZW6+E+22FzwVsXrf
l+D3yHsMjv6qYg7ANCEletDc/JpqBwlE3C+RC7E3lGFyP9TGWymUhNyvlTGBCUsnzP6UDJuDWVzQ
tCtd/LxB+Xazv/ZXyO6ClMf8z5s0ogBic6LUVSbKkWXXuWaob8wMYug2O2gTQ0gVJAxjn18vrVpU
tqGHaI8hEw6PCvyVkj/Lp76YnA22q0XoV2V1oFH13x20iZAUndPCh+o1TarWWHDq9tmjO43s9axl
fFRza9Ri5H/2yDpw4SCx+Ia5geFRwS52mHBLwnhrKh6GH4xmMxEUW55hjUsUk9sjCOVbWR/aINCw
2r3nch8xO3snTM1F78gp0+KvVKl8oxNCtR+5eGO3VrDWX+B3YgdsUngfu+xP7Bu/R2d2N9yJWjE8
dzEsWQPK2zgKNaS4xdFo8kR9fdtgR0ZPGMeRvPKWNcO9HfSa8c4vVgvvstkZR7Z04Kl4VD4Tw9ry
4tq32Ox3COqZBVxDhRI8cJBgY/URSs2MetzgGWHm5aMnmVB/8kPe641LtroUW6APZ8DhyFtdkmUI
p5wT1r+wVQV/be2KntxWrqgGC2XltqNXL/McwaJ4a25QFvXJ2iTeS2WlKwwQYPvz70P3NZJMhKYD
5igDJkMvubdPR0h0CEepAkRZr9aS6lNZKVj8HyOM9KgoK/tBrb3tVw2Hh9ejKUdeY9aUOMPKy3My
xofKBbRQxQmZ9n8nFkDbrdujm4v+60fm87F3Y6AF1Ddjv0wI+TLUyLiNY33g1/yGVdqkPOqAeX8/
SvLZ3IVhIdkAnYzbCZ6xznnMyUEq+s3231y20PKqb7KldIGLcUn5hAeFw7cj2Ui1rdJclIsrumvI
lLM5I7/B4vDW9/Zojn8HvENRDUf1vMg58qptM1rHx5ToxCy9Oo/P6paazktxsWIsph7R7LbN9TDU
m1kHsIKejs4Ch04Hg2rCf+iCR13PQZfB9zYbCYEMz6Fk3NOQK5nuHBrOMPh0clnm4OzzezZSAt0b
zVK+TXNwdi2pzMrezO/2VX/vQr5iZZsu7x4QgGz+dIwsRL53ygVtDfOhIXuw3PJMKa/aAHCiLuSM
BzJHjHzgTZwheV+UnLTYb1PJcUOSZqhHd1mFGSD+vRzjfuUq22CTEPX+6qyqs6EswPGUDCJpKJ+B
nzmBKOGXocS2E00YH96IJyRzqg/LO1aynhaSzVkLw6v3dhqA/Pyr352fEVGwyDR9ESb4p9/aDiev
F4nNHCqlUEvgfe31jyeutvSwyFiP1U0nF3sWXSL3ys/zVjjlXu4kGGBpwAJDQBjVPfUaw4mWS2j/
+/UsOGl52hYtrj2LRztx6zp0tcRXxkyyiOBuF4YWOqG/UKUOBda66I5Eiy/YKjOEl4WGOjjejgs6
ed07jnYhUXqBLWp7bemeEVKFJJETe4e3ZCLqDkgHJEekMivTQxpZxHTu1ZrQziGNe5M8JrPQDDiQ
crtvknPmnsKOW1TjCBgYMFTujHoIiajZbRlBJkMa9qUvtX4nEmksjg7fTxmNcuziYhX9mUyXhHWm
z6LiO00giBqutd70gS3PiyHtNBz34tOvnBIXVMzHkdqBnIZQRlCX9el5B7dXHktHcFaaVC7qyKXs
3PQdcWUaDYJpMT4+YefgRmOL6beahNL4n1kusIlsRBtxFfzMCqbqjFBG4xhtpBgi9Q5t2N2uDlM8
/a1vdpWUubdzBT2hRJol/YFmjKTH74IIbziX24s3pR40Tt3F0bxgufQ/tCQgCzO7Fg6Yd0407XF/
PmWk1F80zhwj8VGr4JV9pihFVEmAZr0af/hAE++GiwlXdZcFsRyphNjVYS8Ev12GdNjTJk5eZFfH
22yytaQGG9BqFyJqzn9fLuqc4hyPnFVeoN+B/rOPm/ZEP/M8Z95qll6txVsYLbbRkJ/gyNtCn4KX
ees/QeY6C9GSOVzTtp9jiQ0qkdhTZjiaOQam1aFMz4OpRtNuBGKQyDXAb2ATcPNUsoq1XXifq6Wf
EG19yXcf837jQ4qw0S5+DfF9aOIW0I9OmXhoJ52dBo0RrAYdjOv2/1HzFj2sAzo6cAqBbdbZ6n0B
cfJIFylXLyW7EDzJJpzOAeIJ30+3RaI7zGCcOHq7yQg6ushx7qtFlmiw4lJzqdKgu3BjoZbsdIuD
SbWEWrsObczgugI5VNOB6c5vrJTpOzUiRUbNcImdRDiVNLqwwz7fwWIE2W22dATUsqJ5FQYfUp1E
eMa/FWH/pF45oBSXaOUDNbxmkh/5TXFBkfyYAW9ImB4dYEvSDh+ISne/9R0qVMOgNoTRuhjy2Rr8
q8dAPlulMDOTdtsZ/LS9c1NNTw88pqFktSVtoEOo7KZ9iRV3gwh3oE9mKaLRlpt2evmA5Ako+kxd
qd8s5tbeeoeccKr4txAWLDcKuOgCiqLzWjBWUcg9YWX+f59sB+L3kQkNihDsJWRGd55ImsI6+zQ/
KIA8KMae6MBM1KL45o4pxZKmOZuYkz69nGM4qUaZWXRcBKGjgwebzrINggggET29HDOeUIBlocV5
Vx6hnU3wSlIXZrLgxPGJsfwbH5iamrNf7yL0GGO9RSmSKHZQP5Y+wFIwAb2PN/rapzpD8Ldkg1uO
kE5KR8uH0+BvUy8okipfa+iX4s2KrTSbuSGwJWyYM+zu+U25dyTnjAm5s7XWzhW+y2/rAsAcfyC0
dtzw4wPe+qvISszBjEJhzv2Z1hQrf8fmLWT4JxEvmdfahExg8eoHYPanlDYKKpNKX0aJOVPZstJp
jg2Ca2T11tlkYh6NLK9/04W7yYfHfpcokjNRm/nm+3AHh+QRd7fvaJpIPpSPDt344fVjiFocL8ZC
VE0kZgTz0ZbkMaxdXXp1di1p5fGuZ18SLjIzvfzmjhHVS+zccNJvSUGE+N8ZNjtscf1rAO4umVkv
iXSV0cxkCxb08WKeKI46dexd5yAQHziV2BuavtXo7zx3d4KqrxGnELX5+UzohUaPkyQScQ8hMPiW
lY0fWK0fc2IGMKUehfJZVz0G41i6lKNovH/Rwyp3BZgZ+sVXHMfHBtXRtjmqXsk5Kouqeou7LISs
iBKO/lwXyxTaSk9PZgLxk7Lwg9gjS4LzIKllz40xRZm9ApFYsZ4hb6NexUb4vUAp+cs5qQPDiLxJ
3qOrr2hLI52WGldE3Blni5Oz9WmHAjPY4sCTX53gS6DC014QXiGJncSIp+m3tXrbBRGKzt7iLpvq
Pph1vMFEDi0hqmfaGQh5f2O/nq/flUNqUyAmzv3Puen/da2ThU3nQ2XfPeGbBOdmMi52wOLCHJYr
qyE9gIZ8bC6i1BMKWvYUNh4GySYkYvkBDPpJHnlrjoxoqBu09RVrAAObzubepzSXo8pG0fl1DGdy
HdvM6K0BUGwZUZjuiKpChxDSti+u3GlMwhUnVQlYMhguED+yCW9yLdSfM3vqZ3JQafeSsUKz0s0x
l915E/rbGsqQhVu+OQGxjAJUoz4UcB78abtahIgR9fQU4Fs1SD90Bg/TBoYIwKaW+7mWzp6RK5sH
jKHonLVMPRvKP126JUWdQfLxqLQYcPLcaLoA/xb2RqxF2Zu8t0BtYrIg8hLecGPfn87vjxD5fh57
8uJAj5FFX+yKXlWsGKFAaeFaAvXRhcQlQksrn8Jfj9pbVZxIV/oRI7D132XZ57lI4cbL/bb1QDtU
ucyZ33t3ftjgcW7p+T9vEAsbEU6yDnjfC7UlVSGmhCimviJ+6FZBonWFD6oh/twLeUFVztKnswAE
XheWZghGXc1FO9oyJ+arvb6RJwj77FJTIhMHpyWNIb7SN5CB8v51hOvW7Yn5KJXmrJcfWC/27Stg
dORY8ZuSsruXsx/o2zzm5xvH9kA2XA0npyAgw5SsG9TchmDKBTMF5uwi6SZzBOvt+b/VDePLRch2
C1zaUP1lHi0A0BAiVIV8zyvaJIwCrArMK9XWmmEW8ru2q+IYT2ac8RC4tP7a9eDaCIIfYu1FIqLx
IcwfeZonUMKq78C4Pk8mBxbIGGB0n8AmKHhPAwgr7iqk28cjB7zkEVC5VCjMymnFN35Yyx0hP1+A
VQg2t6MNJ4bUQAcRFcVLy7UMevn76enCkI81Cqmh17CE4F3zLjw9zio4XsuS/k2SknfnprTxqY4Z
D8CvP4dI78V9leMAHJxP8atdrZl7CKkgAZVKPykChA+wvO+5jZASUQEHJyTf0GxZZ/Uw9JywR5CL
7W5d3S4iQSXgfLAzdeDEcwtxK148anh4Rq62xwX5E2xXHKOps4FeOTW8fC7rPXCRpIiHtN3+ZraI
Ex1+jLJMwkvPKnDc9aZnnuMkMJ53mCoJt4irFKJEQGezYGGh8W1SI8+uvgmSb2JrYH1he18wdnKL
UTSsdtZ+cgVvcFVmS2gnkZhse4h/km/450L/Izlnj3fB8tMKLraCyDvyvbtlsOS/Wmp5i6Bd1EQy
Vb+ubzp5VR8XDE0a44HvERdI/3SRPb4nBJD6YJ2W1CPKDpNP9FafiVPG+CC3zrhTiWpgupp4r7H3
1h1CSDUSd39tztQcyZMsMDUFzHWYW02IDtFZnBSIJHKQhToVVVSmhmbWPCizIi9edykzq5ABdpV0
6kR3DorPGOfkL3ZAka7Ot39FhVX8BQDUwiUo9Tt47WRVNdiQJ/UHJ2fQh7/2miu7rpPJu3m6h0fw
puW6vI/GN+eL3nk4W5LOmSnT4cnON3n1Ev9bZGySlAEN7vzDSNjBKoc6z88A+KgOnqqyt65MqPr2
NEYfuT8Zq8Cd2lrCqWOFUPSVOaTal8FbLaBlAHBiwXDJ1RwiInm1j4l1qJpBtt+5ydtKoCMc5UAb
ziA3TUGT9PxcqLt6ZzXaR5BVK6zzBRYw5r9o4GXQQRZiUvqUkqMhFj2TB3PlhDOzb8m0gdF7/fGw
rYf0d10KaY40q4Bku2uPZtMGi8Trh82SFLgJO1+xXmM7K/WgpuN6TUx8A3fFJ4IgUqOd7weJMOAP
b2cqSM10wT9rtMnhEsKDBDRKKvniY7DHUYOUQqKSuVgdT7coyBEdELs9z/Hr3YEl7Hw8BY2spMNM
ib9Z2a8pm8M/Cc53mlKIyYJPOUYxNhY96ysVTwBp4ULSu7mK65xDMRlS8rm9SGAsf/9AlgiqLNGc
18RxU5K/ztpM0T76PJpvEUgV66TANCEuobpbS3cY/vVk3JBlUwGaF16HLdaUpsYyPjpy1lUyl5CX
jemb4ryxX7sMQL9M5A3hfHiAOtXJBibh2uS7+kBXlX+AOuMwCcp9e3ZFtGJFP0fn1b1EARLvoiZF
YiDxmeOAdu75nrPZJGnofCR0ca+cfRV5jwR1U9KJjwd7jGYaDP7NLzzBfg7yAmFsYPd03QB6Vr5y
BiXgjI5ub2nYbbaAmppN70EAuPuPH0ZD6Epe7nNx0kotgqJ8A3w9SsunU/h9TIH6nq0yvc0En9If
tlUeg8p5CdmCUK8Sz7WR+IBNJyhsv90baWVfL7TsUxfr5cFJJbk6dPwyf5evU9jyM6kovAuIngGb
dRhCrXD22IZ+YuoQxAlfqKv2oMO+aITvFCyWYYAA1UCpLE/ze7+EGolApFuhfWn09gKhHAsVJTvh
geNM9WHweOfO3ic1u6Ab28ee7tZLAEB0I5jal9kel2/6gtI4XfcAQyZvvsiqEPcvZk4xMvpu71mw
wTl/TdEziwPuqQZGzFGjekutnclGw6i49KYxDaUm1wtOXpVnOLAtejnGnrQXVstgXl5PfZ+72jak
G5w4e82/EvCKgO7rbESZltl/gCZ+ARTZEvGk/nkPJQl95NjoFxVGPBv5M9Ob3f7YJnFK5AXoBULW
Pqi0pm7+lCOMsvnqTVPR06wQ2twdr2/YRcaWlHZlSfG2mYkByviXSjTvlkvXATqkjU+FLZJK1I9C
MfC9D1a8FtH3EOk2DTiu5pIPLn2C8V6+w/Mv0HwChU/0bOmU6Yg/unHjmK5D0dPahLbSNpV6n0ui
Pto7ByEeo6Bq7A1N1X3s4TtmnncWe7BQuCp500V/ViOc7gMJLT/Z+nakLDiCjzTYfrNEv0mqppRj
nmvUPW0cm2JIFDOj1rOe4inQln3jZo7XRJTr7WvbskDbkVG74LFNGiyIRzCYiQ/sWzrxKFpy8Ns5
DP0CTi+2FV/K1WAmhfhhmoYKaAGkeWQ6tKkyb6IWzojqfONlTZNuaN8Jss5QOiuoqTDOLzx9altw
feDfygMI6POP7K/lWRhqM5uDeRv1WWedMaslg0zCezYRInWrIYgmu/0/KQlqoXY2L+kQhQzwIgPR
0GIyIre3yYBsY/BRvDAcuGdAsETurZTATRqTS1kcYoYr6s8rgQD/7bWpLqxbRidQH6YoUKxo9yQ3
2VwZ4/GpPIWkAMvHqouN6Z20+UTysYwVnQJnEMW2i1rVfzWhXPw/MbuRfUsKyT7G20hjEqO49KWP
i2vHPeUnvCZrx6d6KntApk9RabZ+IAu8+ZKhpB6i6k64vhkmLoZHWWxSP2tnTfOV2WW0Ld88lpzN
3lPJE5jDueh5y+dVuToHmaUSPExFCf/pQDODvr+nFBprPrLiRpEjXVROlKJ96Z0Ub3Te08/s2fn0
ZnmvwD3/rNy1y0lHgpU+7VkjZjkvFpZjhINLK+Nmruao9q9yfXqydCaulH4ER+fq6166W6eMHIEN
tjInRsMpiCKPM4lTB4WWDK0w4E2skc8eiNks7vaGr1+Fw3KItxnKoyOB8lxEWu65s1Ptc6h/77iP
9bb8QwSbR3DVWUTGQDGj0B3HX+FcHaEil4i7sCWJdkI2kW5O5Whq99DvT65M7LsTZ2z9skgkCWIH
g7MhugvsGN7ItZ+H4hRjZM7YerhmKLVp2Uar2ralT56ZQ21a5o26wbv/VzPBTrBfujhEXqs8mQK/
LTvpAr2jA+tzipCo+aiJ4IxISgv/iApiS8/OpGbteiGn93zAiqREd+7Db2dYrRo0ICTNKFzT6588
Wn9BS+mA1RG1vmLwxFOsvXV5/VTnYhpt5kd7fWbTuBB46xOoL3vpdfxZ6a/+DkqC4JZBk3G5e1d3
rX7o0Dtj0nsNUWmYezYSC+TCrarb5pdQtZ9Mjc3LizwzNBIl6yyu6KjXTXN97Ofctwbg3qhQ9t7r
TdGqu71NkRPBF923oypdpAt9cBr/IPv1U/SXb92sATwSyezVCF0VDHKEjdQV/6eZCI1yc02YPiew
RNwqoO3H4GeumRWW1s1tIY/dCG3cA5dFNKDe3xHLZtB7ajr7ll/EeZQ2XEP8SU9Sx0s8bhhV2KeM
AeSQ0dXuqwv+gJnj933NyDLYm3fG7624JAN47GGhZl15qq/4fazVvNperlQQMPqx0bNQ9pbn93ZL
WKtajDT32jztbHHirJhiXG6dJQRO45lEzcKaLbgJtQdp5j9ycN/dyxyBgO2+H0ybpHKwW8UAUS6k
R5svcmiHTjn+nT0yN5qGPv186e2f1NkmoAhj86t7JOwLN9Os0sAqWN6P6bqFKX2i+hcq337M1lsZ
vdRkmakT5ah4/zB5cRBjc+DNNH/gQ4MUmVxqg6ZN4c9Ouxv98F594kWnMn+ZSslHf6uulaYJ+io6
yTLZ9mnQMW35Ve15TC8w7ZoLkRUTllG2/gQCpeFN767oVKkqVAbb5B+jqTvByKzBSLPZEFhOsNBS
p4L+LIZA3cQvf/Iq8H2nutCSXCl+Q1CGm1QoLgMrNjKCL4mAZvPK2TC3Ge/VVuAAU6gM6PQfxM5l
8Ok02oaJj5ymvjYv2J5DBLGIIlx4eziJ/Ok5/qV1kwQzRkC/XZdQikW27k2eRCKQtJwmX3qVxCb7
qZOXExK+XGo2JFhl0KlbN0GejRP7FGA4HWPoAm2h9FOH4x2ISj2zJxdFYKSlA4NvPmm/Ptt2/Wu/
Pbc3Mjm5tobjZvYoEWVbarr4B+NGSIWhDmRW77L/BS1npY5F7Knixh2h35IpIyCN/E1Uly9e5TwZ
OIr59pGOlDxZA843oTW1MHzLKOKfygO2G2IaAtUjzwXk3LxGteUlDEaiFOw4wfJEdFKAxW2C4ueg
accq2KmG59SBssNxOD4hlD6hBAsFG87g5uVTKlNjtXzmElkVl1TKEMWreI9vXODfOybJAvghhGPe
JQqE9W63s2eGgCmQaheo+xdVAMMHZIhh5vnRnaDY6XUq0WJ8fbxGGkN6C2u7i9Ni5FgCorKUJBIt
OWJLj++6Deof2EjDQsb0gQIx6s+YdVlVdftHH4v0TPvFjGjXJ5eHGRGGQEkHxFOI/YI/Deyh2+md
Ss91zAXlWCbX4HwszvKegvXB/J9LnMwTJTfcUw5ireASYzezyI5EMYpXaNMUHIeRYheZ9bz+IAdn
qqP03dWU2jYvy08wlbQYtsL5RxmsY/pJbH0OFDBMjsQBV9yd6+05u+uaqUrLhHHd38iCsWQzCVUT
vYrZ/bW+VOx4RbHcFd561piawYNeVKG3pACe5AnJ99JwlQQLPSHlUIXOcfDEI8RDI2aSjS8opmE3
8/hYuYQtpsG38tJlTAlfiRkvSUnjF0zGhDGPxQ5eamPdkM41I4+5JdDBDSOCySaPsY7ySZlm1i1x
w4VsIb5IhRSHMFM3CgT77k7DAX5DS2/jCmthbCURMbYAOPssc9fikUeL1ORLZfLLtKeKpTS769Bb
MROXXaSbVmYLhY9+wZ1irxi7fWMjSGEM69CAS9XZUYUi9WvWrAZRkXn8ceXa6qwPLkFwZ5rI4eFh
bM145SjQncuLgy2ee7FxL3KKUEeDfxo3jPn8Z5sk+T5/L/PNuYpvE3D5NjhFFoRTjWf4OdIkZ+Ef
HcWQqZk8+ukloEONWz3wUdsV0TYURCKqjnrirWgWLlJS1m4PVNIWREgpvGIrfYLPudp+I2HQ6e2s
TScBHlZdl87P2dMRJmPey5BNnOaJOTLDdW4cvL6J
`protect end_protected
