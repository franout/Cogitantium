`ifndef __PRECISION_DEF_VH
`define __PRECISION_DEF_VH


`define  LOG_ALLOWED_PRECISIONS 4 //LOG 2 of total allowed precions (9) 

// integer
`define INT4 4'h0
`define INT8 4'h1
`define INT16 4'h3
`define INT32 4'h7
`define INT64 4'hf
//FLOATING POINT
//TODO CHANGE 
/*
`define FP16 4'h5
`define BFPP16 4'h6
`define FP32 4'h7
`define FP64 4'h8
*/
`define VIVADO_MAC 1


`endif