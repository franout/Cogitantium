// Register NVDLA_CSC_S_STATUS_0
#define NVDLA_CSC_S_STATUS_0					32'h4000
#define NVDLA_CSC_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CSC_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CSC_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CSC_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CSC_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CSC_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CSC_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CSC_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CSC_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CSC_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CSC_S_POINTER_0
#define NVDLA_CSC_S_POINTER_0					32'h4004
#define NVDLA_CSC_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CSC_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CSC_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CSC_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CSC_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CSC_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CSC_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CSC_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CSC_D_OP_ENABLE_0
#define NVDLA_CSC_D_OP_ENABLE_0					32'h4008
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CSC_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CSC_D_MISC_CFG_0
#define NVDLA_CSC_D_MISC_CFG_0					32'h400c
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_RANGE			9:8
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_SIZE				2
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_INT8			2'h0
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_INT16			2'h1
#define NVDLA_CSC_D_MISC_CFG_0_IN_PRECISION_FP16			2'h2
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CSC_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_RANGE			16:16
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_DATA_REUSE_ENABLE			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_RANGE			20:20
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_WEIGHT_REUSE_ENABLE			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_RANGE			24:24
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_DATA_RLS_ENABLE			1'h1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_RANGE			28:28
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_SIZE				1
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_DISABLE			1'h0
#define NVDLA_CSC_D_MISC_CFG_0_SKIP_WEIGHT_RLS_ENABLE			1'h1


// Register NVDLA_CSC_D_DATAIN_FORMAT_0
#define NVDLA_CSC_D_DATAIN_FORMAT_0					32'h4010
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_RANGE			0:0
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_SIZE				1
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_FEATURE			1'h0
#define NVDLA_CSC_D_DATAIN_FORMAT_0_DATAIN_FORMAT_PIXEL			1'h1


// Register NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0					32'h4014
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_WIDTH_EXT_RANGE			12:0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_WIDTH_EXT_SIZE				13
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_HEIGHT_EXT_RANGE			28:16
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_0_0_DATAIN_HEIGHT_EXT_SIZE				13


// Register NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0					32'h4018
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0_DATAIN_CHANNEL_EXT_RANGE			12:0
#define NVDLA_CSC_D_DATAIN_SIZE_EXT_1_0_DATAIN_CHANNEL_EXT_SIZE				13


// Register NVDLA_CSC_D_BATCH_NUMBER_0
#define NVDLA_CSC_D_BATCH_NUMBER_0					32'h401c
#define NVDLA_CSC_D_BATCH_NUMBER_0_BATCHES_RANGE			4:0
#define NVDLA_CSC_D_BATCH_NUMBER_0_BATCHES_SIZE				5


// Register NVDLA_CSC_D_POST_Y_EXTENSION_0
#define NVDLA_CSC_D_POST_Y_EXTENSION_0					32'h4020
#define NVDLA_CSC_D_POST_Y_EXTENSION_0_Y_EXTENSION_RANGE			1:0
#define NVDLA_CSC_D_POST_Y_EXTENSION_0_Y_EXTENSION_SIZE				2


// Register NVDLA_CSC_D_ENTRY_PER_SLICE_0
#define NVDLA_CSC_D_ENTRY_PER_SLICE_0					32'h4024
#define NVDLA_CSC_D_ENTRY_PER_SLICE_0_ENTRIES_RANGE			13:0
#define NVDLA_CSC_D_ENTRY_PER_SLICE_0_ENTRIES_SIZE				14


// Register NVDLA_CSC_D_WEIGHT_FORMAT_0
#define NVDLA_CSC_D_WEIGHT_FORMAT_0					32'h4028
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_RANGE			0:0
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_SIZE				1
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_UNCOMPRESSED			1'h0
#define NVDLA_CSC_D_WEIGHT_FORMAT_0_WEIGHT_FORMAT_COMPRESSED			1'h1


// Register NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0					32'h402c
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_WIDTH_EXT_RANGE			4:0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_WIDTH_EXT_SIZE				5
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_HEIGHT_EXT_RANGE			20:16
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_0_0_WEIGHT_HEIGHT_EXT_SIZE				5


// Register NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0					32'h4030
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_CHANNEL_EXT_RANGE			12:0
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_CHANNEL_EXT_SIZE				13
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_KERNEL_RANGE			28:16
#define NVDLA_CSC_D_WEIGHT_SIZE_EXT_1_0_WEIGHT_KERNEL_SIZE				13


// Register NVDLA_CSC_D_WEIGHT_BYTES_0
#define NVDLA_CSC_D_WEIGHT_BYTES_0					32'h4034
#define NVDLA_CSC_D_WEIGHT_BYTES_0_WEIGHT_BYTES_RANGE			31:0
#define NVDLA_CSC_D_WEIGHT_BYTES_0_WEIGHT_BYTES_SIZE				32


// Register NVDLA_CSC_D_WMB_BYTES_0
#define NVDLA_CSC_D_WMB_BYTES_0					32'h4038
#define NVDLA_CSC_D_WMB_BYTES_0_WMB_BYTES_RANGE			27:0
#define NVDLA_CSC_D_WMB_BYTES_0_WMB_BYTES_SIZE				28


// Register NVDLA_CSC_D_DATAOUT_SIZE_0_0
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0					32'h403c
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_RANGE			12:0
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_WIDTH_SIZE				13
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_RANGE			28:16
#define NVDLA_CSC_D_DATAOUT_SIZE_0_0_DATAOUT_HEIGHT_SIZE				13


// Register NVDLA_CSC_D_DATAOUT_SIZE_1_0
#define NVDLA_CSC_D_DATAOUT_SIZE_1_0					32'h4040
#define NVDLA_CSC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_RANGE			12:0
#define NVDLA_CSC_D_DATAOUT_SIZE_1_0_DATAOUT_CHANNEL_SIZE				13


// Register NVDLA_CSC_D_ATOMICS_0
#define NVDLA_CSC_D_ATOMICS_0					32'h4044
#define NVDLA_CSC_D_ATOMICS_0_ATOMICS_RANGE			20:0
#define NVDLA_CSC_D_ATOMICS_0_ATOMICS_SIZE				21


// Register NVDLA_CSC_D_RELEASE_0
#define NVDLA_CSC_D_RELEASE_0					32'h4048
#define NVDLA_CSC_D_RELEASE_0_RLS_SLICES_RANGE			11:0
#define NVDLA_CSC_D_RELEASE_0_RLS_SLICES_SIZE				12


// Register NVDLA_CSC_D_CONV_STRIDE_EXT_0
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0					32'h404c
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_X_STRIDE_EXT_RANGE			2:0
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_X_STRIDE_EXT_SIZE				3
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_Y_STRIDE_EXT_RANGE			18:16
#define NVDLA_CSC_D_CONV_STRIDE_EXT_0_CONV_Y_STRIDE_EXT_SIZE				3


// Register NVDLA_CSC_D_DILATION_EXT_0
#define NVDLA_CSC_D_DILATION_EXT_0					32'h4050
#define NVDLA_CSC_D_DILATION_EXT_0_X_DILATION_EXT_RANGE			4:0
#define NVDLA_CSC_D_DILATION_EXT_0_X_DILATION_EXT_SIZE				5
#define NVDLA_CSC_D_DILATION_EXT_0_Y_DILATION_EXT_RANGE			20:16
#define NVDLA_CSC_D_DILATION_EXT_0_Y_DILATION_EXT_SIZE				5


// Register NVDLA_CSC_D_ZERO_PADDING_0
#define NVDLA_CSC_D_ZERO_PADDING_0					32'h4054
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_LEFT_RANGE			4:0
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_LEFT_SIZE				5
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_TOP_RANGE			20:16
#define NVDLA_CSC_D_ZERO_PADDING_0_PAD_TOP_SIZE				5


// Register NVDLA_CSC_D_ZERO_PADDING_VALUE_0
#define NVDLA_CSC_D_ZERO_PADDING_VALUE_0					32'h4058
#define NVDLA_CSC_D_ZERO_PADDING_VALUE_0_PAD_VALUE_RANGE			15:0
#define NVDLA_CSC_D_ZERO_PADDING_VALUE_0_PAD_VALUE_SIZE				16


// Register NVDLA_CSC_D_BANK_0
#define NVDLA_CSC_D_BANK_0					32'h405c
#define NVDLA_CSC_D_BANK_0_DATA_BANK_RANGE			4:0
#define NVDLA_CSC_D_BANK_0_DATA_BANK_SIZE				5
#define NVDLA_CSC_D_BANK_0_WEIGHT_BANK_RANGE			20:16
#define NVDLA_CSC_D_BANK_0_WEIGHT_BANK_SIZE				5


// Register NVDLA_CSC_D_PRA_CFG_0
#define NVDLA_CSC_D_PRA_CFG_0					32'h4060
#define NVDLA_CSC_D_PRA_CFG_0_PRA_TRUNCATE_RANGE			1:0
#define NVDLA_CSC_D_PRA_CFG_0_PRA_TRUNCATE_SIZE				2


// Register NVDLA_CSC_D_CYA_0
#define NVDLA_CSC_D_CYA_0					32'h4064
#define NVDLA_CSC_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_CSC_D_CYA_0_CYA_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_CSC	32'h4000
