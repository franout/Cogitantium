// Register NVDLA_CFGROM_CFGROM_HW_VERSION_0
#define NVDLA_CFGROM_CFGROM_HW_VERSION_0					32'h0
#define NVDLA_CFGROM_CFGROM_HW_VERSION_0_HW_VERSION_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_HW_VERSION_0_HW_VERSION_SIZE				32


// Register NVDLA_CFGROM_CFGROM_GLB_DESC_0
#define NVDLA_CFGROM_CFGROM_GLB_DESC_0					32'h4
#define NVDLA_CFGROM_CFGROM_GLB_DESC_0_GLB_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_GLB_DESC_0_GLB_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_DESC_0
#define NVDLA_CFGROM_CFGROM_CIF_DESC_0					32'h8
#define NVDLA_CFGROM_CFGROM_CIF_DESC_0_CIF_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_DESC_0_CIF_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0					32'hc
#define NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0_CIF_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_INCOMPAT_0_CIF_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0					32'h10
#define NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0_CIF_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_CAP_COMPAT_0_CIF_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0					32'h14
#define NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0_CIF_BASE_WIDTH_RANGE			7:0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_WIDTH_0_CIF_BASE_WIDTH_SIZE				8


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0					32'h18
#define NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0_CIF_BASE_LATENCY_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_LATENCY_0_CIF_BASE_LATENCY_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0					32'h1c
#define NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0_BASE_BURST_LENGTH_MAX_RANGE			31:5
#define NVDLA_CFGROM_CFGROM_CIF_BASE_BURST_LENGTH_MAX_0_BASE_BURST_LENGTH_MAX_SIZE				27


// Register NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0					32'h20
#define NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0_CIF_BASE_MEM_ADDR_WIDTH_RANGE			31:5
#define NVDLA_CFGROM_CFGROM_CIF_BASE_MEM_ADDR_WIDTH_0_CIF_BASE_MEM_ADDR_WIDTH_SIZE				27


// Register NVDLA_CFGROM_CFGROM_CDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_CDMA_DESC_0					32'h24
#define NVDLA_CFGROM_CFGROM_CDMA_DESC_0_CDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_DESC_0_CDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0					32'h28
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0_CDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_INCOMPAT_0_CDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0					32'h2c
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0_CDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_CAP_COMPAT_0_CDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0					32'h30
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0_CDMA_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_FEATURE_TYPES_0_CDMA_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0					32'h34
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0_CDMA_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_WEIGHT_TYPES_0_CDMA_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0					32'h38
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0_CDMA_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_C_0_CDMA_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0					32'h3c
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0_CDMA_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_K_0_CDMA_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0					32'h40
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0_CDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_ATOMIC_M_0_CDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0					32'h44
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0_CDMA_BASE_CBUF_BANK_NUM_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_NUM_0_CDMA_BASE_CBUF_BANK_NUM_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0					32'h48
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0_CDMA_BASE_CBUF_BANK_WIDTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_WIDTH_0_CDMA_BASE_CBUF_BANK_WIDTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0					32'h4c
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0_CDMA_BASE_CBUF_BANK_DEPTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_BASE_CBUF_BANK_DEPTH_0_CDMA_BASE_CBUF_BANK_DEPTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0					32'h50
#define NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0_CDMA_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_MULTI_BATCH_MAX_0_CDMA_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0					32'h54
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0_CDMA_IMAGE_IN_FORMATS_PACKED_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_PACKED_0_CDMA_IMAGE_IN_FORMATS_PACKED_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0					32'h58
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0_CDMA_IMAGE_IN_FORMATS_SEMI_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDMA_IMAGE_IN_FORMATS_SEMI_0_CDMA_IMAGE_IN_FORMATS_SEMI_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_DESC_0
#define NVDLA_CFGROM_CFGROM_CBUF_DESC_0					32'h5c
#define NVDLA_CFGROM_CFGROM_CBUF_DESC_0_CBUF_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_DESC_0_CBUF_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0					32'h60
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0_CBUF_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_INCOMPAT_0_CBUF_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0					32'h64
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0_CBUF_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_CAP_COMPAT_0_CBUF_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0					32'h68
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0_CBUF_BASE_CBUF_BANK_NUM_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_NUM_0_CBUF_BASE_CBUF_BANK_NUM_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0					32'h6c
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0_CBUF_BASE_CBUF_BANK_WIDTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_WIDTH_0_CBUF_BASE_CBUF_BANK_WIDTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0					32'h70
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0_CBUF_BASE_CBUF_BANK_DEPTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CBUF_BANK_DEPTH_0_CBUF_BASE_CBUF_BANK_DEPTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0					32'h74
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0_CBUF_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CBUF_BASE_CDMA_ID_0_CBUF_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_DESC_0
#define NVDLA_CFGROM_CFGROM_CSC_DESC_0					32'h78
#define NVDLA_CFGROM_CFGROM_CSC_DESC_0_CSC_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_DESC_0_CSC_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0					32'h7c
#define NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0_CSC_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_INCOMPAT_0_CSC_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0					32'h80
#define NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0_CSC_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_CAP_COMPAT_0_CSC_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0					32'h84
#define NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0_CSC_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_FEATURE_TYPES_0_CSC_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0					32'h88
#define NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0_CSC_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_WEIGHT_TYPES_0_CSC_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0					32'h8c
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0_CSC_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_C_0_CSC_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0					32'h90
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0_CSC_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_K_0_CSC_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0					32'h94
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0_CSC_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_ATOMIC_M_0_CSC_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0					32'h98
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0_CSC_BASE_CBUF_BANK_NUM_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_NUM_0_CSC_BASE_CBUF_BANK_NUM_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0					32'h9c
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0_CSC_BASE_CBUF_BANK_WIDTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_WIDTH_0_CSC_BASE_CBUF_BANK_WIDTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0					32'ha0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0_CSC_BASE_CBUF_BANK_DEPTH_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CBUF_BANK_DEPTH_0_CSC_BASE_CBUF_BANK_DEPTH_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0					32'ha4
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0_CSC_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_BASE_CDMA_ID_0_CSC_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0					32'ha8
#define NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0_CSC_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CSC_MULTI_BATCH_MAX_0_CSC_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0					32'hac
#define NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0_CMAC_A_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_DESC_0_CMAC_A_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0					32'hb0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0_CMAC_A_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_INCOMPAT_0_CMAC_A_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0					32'hb4
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0_CMAC_A_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_CAP_COMPAT_0_CMAC_A_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0					32'hb8
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0_CMAC_A_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_FEATURE_TYPES_0_CMAC_A_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0					32'hbc
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0_CMAC_A_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_WEIGHT_TYPES_0_CMAC_A_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0					32'hc0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0_CMAC_A_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_C_0_CMAC_A_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0					32'hc4
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0_CMAC_A_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_ATOMIC_K_0_CMAC_A_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0					32'hc8
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0_CMAC_A_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_A_BASE_CDMA_ID_0_CMAC_A_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0					32'hcc
#define NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0_CMAC_B_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_DESC_0_CMAC_B_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0					32'hd0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0_CMAC_B_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_INCOMPAT_0_CMAC_B_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0					32'hd4
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0_CMAC_B_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_CAP_COMPAT_0_CMAC_B_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0					32'hd8
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0_CMAC_B_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_FEATURE_TYPES_0_CMAC_B_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0					32'hdc
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0_CMAC_B_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_WEIGHT_TYPES_0_CMAC_B_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0					32'he0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0_CMAC_B_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_C_0_CMAC_B_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0					32'he4
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0_CMAC_B_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_ATOMIC_K_0_CMAC_B_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0					32'he8
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0_CMAC_B_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CMAC_B_BASE_CDMA_ID_0_CMAC_B_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_DESC_0
#define NVDLA_CFGROM_CFGROM_CACC_DESC_0					32'hec
#define NVDLA_CFGROM_CFGROM_CACC_DESC_0_CACC_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_DESC_0_CACC_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0					32'hf0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0_CACC_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_INCOMPAT_0_CACC_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0					32'hf4
#define NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0_CACC_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_CAP_COMPAT_0_CACC_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0					32'hf8
#define NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0_CACC_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_FEATURE_TYPES_0_CACC_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0					32'hfc
#define NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0_CACC_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_WEIGHT_TYPES_0_CACC_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0					32'h100
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0_CACC_BASE_ATOMIC_C_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_C_0_CACC_BASE_ATOMIC_C_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0					32'h104
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0_CACC_BASE_ATOMIC_K_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_ATOMIC_K_0_CACC_BASE_ATOMIC_K_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0					32'h108
#define NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0_CACC_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_BASE_CDMA_ID_0_CACC_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0					32'h10c
#define NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0_CACC_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CACC_MULTI_BATCH_MAX_0_CACC_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0					32'h110
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0_SDP_RDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_DESC_0_SDP_RDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0					32'h114
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0_SDP_RDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_INCOMPAT_0_SDP_RDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0					32'h118
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0_SDP_RDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_CAP_COMPAT_0_SDP_RDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0					32'h11c
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0_SDP_RDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_ATOMIC_M_0_SDP_RDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0					32'h120
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0_SDP_RDMA_BASE_SDP_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_RDMA_BASE_SDP_ID_0_SDP_RDMA_BASE_SDP_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_DESC_0
#define NVDLA_CFGROM_CFGROM_SDP_DESC_0					32'h124
#define NVDLA_CFGROM_CFGROM_SDP_DESC_0_SDP_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_DESC_0_SDP_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0					32'h128
#define NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0_SDP_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_INCOMPAT_0_SDP_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0					32'h12c
#define NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0_SDP_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_CAP_COMPAT_0_SDP_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0					32'h130
#define NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0_SDP_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_FEATURE_TYPES_0_SDP_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0					32'h134
#define NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0_SDP_BASE_WEIGHT_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_WEIGHT_TYPES_0_SDP_BASE_WEIGHT_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0					32'h138
#define NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0_SDP_BASE_CDMA_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_BASE_CDMA_ID_0_SDP_BASE_CDMA_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0
#define NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0					32'h13c
#define NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0_SDP_MULTI_BATCH_MAX_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_MULTI_BATCH_MAX_0_SDP_MULTI_BATCH_MAX_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0					32'h140
#define NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0_SDP_BS_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_BS_THROUGHPUT_0_SDP_BS_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0					32'h144
#define NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0_SDP_BN_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_BN_THROUGHPUT_0_SDP_BN_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0					32'h148
#define NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0_SDP_EW_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_SDP_EW_THROUGHPUT_0_SDP_EW_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0					32'h14c
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0_PDP_RDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_DESC_0_PDP_RDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0					32'h150
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0_PDP_RDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_INCOMPAT_0_PDP_RDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0					32'h154
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0_PDP_RDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_CAP_COMPAT_0_PDP_RDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0					32'h158
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0_PDP_RDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_ATOMIC_M_0_PDP_RDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0					32'h15c
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0_PDP_RDMA_BASE_PDP_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_RDMA_BASE_PDP_ID_0_PDP_RDMA_BASE_PDP_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_DESC_0
#define NVDLA_CFGROM_CFGROM_PDP_DESC_0					32'h160
#define NVDLA_CFGROM_CFGROM_PDP_DESC_0_PDP_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_DESC_0_PDP_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0					32'h164
#define NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0_PDP_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_INCOMPAT_0_PDP_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0					32'h168
#define NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0_PDP_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_CAP_COMPAT_0_PDP_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0					32'h16c
#define NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0_PDP_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_FEATURE_TYPES_0_PDP_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0					32'h170
#define NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0_PDP_BASE_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_PDP_BASE_THROUGHPUT_0_PDP_BASE_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0					32'h174
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0_CDP_RDMA_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_DESC_0_CDP_RDMA_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0					32'h178
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0_CDP_RDMA_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_INCOMPAT_0_CDP_RDMA_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0					32'h17c
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0_CDP_RDMA_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_CAP_COMPAT_0_CDP_RDMA_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0					32'h180
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0_CDP_RDMA_BASE_ATOMIC_M_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_ATOMIC_M_0_CDP_RDMA_BASE_ATOMIC_M_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0					32'h184
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0_CDP_RDMA_BASE_CDP_ID_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_RDMA_BASE_CDP_ID_0_CDP_RDMA_BASE_CDP_ID_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_DESC_0
#define NVDLA_CFGROM_CFGROM_CDP_DESC_0					32'h188
#define NVDLA_CFGROM_CFGROM_CDP_DESC_0_CDP_DESC_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_DESC_0_CDP_DESC_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0					32'h18c
#define NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0_CDP_CAP_INCOMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_INCOMPAT_0_CDP_CAP_INCOMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0					32'h190
#define NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0_CDP_CAP_COMPAT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_CAP_COMPAT_0_CDP_CAP_COMPAT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0					32'h194
#define NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0_CDP_BASE_FEATURE_TYPES_RANGE			11:0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_FEATURE_TYPES_0_CDP_BASE_FEATURE_TYPES_SIZE				12


// Register NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0					32'h198
#define NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0_CDP_BASE_THROUGHPUT_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_CDP_BASE_THROUGHPUT_0_CDP_BASE_THROUGHPUT_SIZE				32


// Register NVDLA_CFGROM_CFGROM_END_OF_LIST_0
#define NVDLA_CFGROM_CFGROM_END_OF_LIST_0					32'h19c
#define NVDLA_CFGROM_CFGROM_END_OF_LIST_0_END_OF_LIST_RANGE			31:0
#define NVDLA_CFGROM_CFGROM_END_OF_LIST_0_END_OF_LIST_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_CFGROM	32'h0
