// Register NVDLA_GEC_FEATURE_0
#define NVDLA_GEC_FEATURE_0					32'he000
#define NVDLA_GEC_FEATURE_0_NUM_ERR_SLICES_RANGE			5:0
#define NVDLA_GEC_FEATURE_0_NUM_ERR_SLICES_SIZE				6
#define NVDLA_GEC_FEATURE_0_NUM_ERR_RANGE			31:16
#define NVDLA_GEC_FEATURE_0_NUM_ERR_SIZE				16


// Register NVDLA_GEC_SWRESET_0
#define NVDLA_GEC_SWRESET_0					32'he004
#define NVDLA_GEC_SWRESET_0_SWRST_RANGE			0:0
#define NVDLA_GEC_SWRESET_0_SWRST_SIZE				1


// Register NVDLA_GEC_MISSIONERR_TYPE_0
#define NVDLA_GEC_MISSIONERR_TYPE_0					32'he008
#define NVDLA_GEC_MISSIONERR_TYPE_0_CODE_RANGE			5:0
#define NVDLA_GEC_MISSIONERR_TYPE_0_CODE_SIZE				6


// Register NVDLA_GEC_CURRENT_COUNTER_VALUE_0
#define NVDLA_GEC_CURRENT_COUNTER_VALUE_0					32'he00c
#define NVDLA_GEC_CURRENT_COUNTER_VALUE_0_VALUE_RANGE			8:0
#define NVDLA_GEC_CURRENT_COUNTER_VALUE_0_VALUE_SIZE				9


// Register NVDLA_GEC_MISSIONERR_INDEX_0
#define NVDLA_GEC_MISSIONERR_INDEX_0					32'he014
#define NVDLA_GEC_MISSIONERR_INDEX_0_IDX_RANGE			6:0
#define NVDLA_GEC_MISSIONERR_INDEX_0_IDX_SIZE				7


// Register NVDLA_GEC_CORRECTABLE_THRESHOLD_0
#define NVDLA_GEC_CORRECTABLE_THRESHOLD_0					32'he018
#define NVDLA_GEC_CORRECTABLE_THRESHOLD_0_COUNT_RANGE			7:0
#define NVDLA_GEC_CORRECTABLE_THRESHOLD_0_COUNT_SIZE				8


// Register NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0					32'he01c
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_RANGE			7:0
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_SIZE				8
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_LOCK			8'h0
#define NVDLA_GEC_MISSIONERR_INJECT_UNLOCK_0_VALUE_UNLOCK			8'he1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0					32'he030
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR0_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR1_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR2_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR3_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR4_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR5_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR6_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR7_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR8_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR9_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR10_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR11_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR12_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR13_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR14_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR15_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR16_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR17_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR18_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR19_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR20_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR21_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR22_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR23_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR24_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR25_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR26_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR27_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR28_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR29_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR30_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_ENABLE_0_ERR31_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0					32'he034
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR0_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR1_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR2_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR3_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR4_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR5_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR6_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR7_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR8_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR9_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR10_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR11_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR12_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR13_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR14_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR15_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR16_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR17_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR18_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR19_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR20_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR21_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR22_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR23_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR24_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR25_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR26_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR27_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR28_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR29_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR30_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_FORCE_0_ERR31_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0					32'he038
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_STATUS_0_ERR31_SIZE				1


// Register NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0					32'he03c
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR0_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR1_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR2_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR3_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR4_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR5_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR6_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR7_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR8_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR15_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR16_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR17_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR18_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR19_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR20_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR21_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR22_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR23_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR24_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR25_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR26_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR27_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR28_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR29_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR30_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_MISSIONERR_INJECT_0_ERR31_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0					32'he040
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR0_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR1_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR2_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR3_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR4_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR5_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR6_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR7_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR8_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR9_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR10_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR11_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR12_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR13_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR14_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR15_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR16_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR17_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR18_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR19_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR20_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR21_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR22_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR23_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR24_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR25_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR26_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR27_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR28_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR29_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR30_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_ENABLE_0_ERR31_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0					32'he044
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR0_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR1_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR2_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR3_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR4_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR5_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR6_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR7_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR8_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR9_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR10_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR11_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR12_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR13_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR14_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR15_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR16_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR17_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR18_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR19_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR20_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR21_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR22_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR23_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR24_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR25_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR26_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR27_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR28_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR29_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR30_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_FORCE_0_ERR31_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0					32'he048
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_LATENTERR_STATUS_0_ERR31_SIZE				1


// Register NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0					32'he050
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_RANGE			0:0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR0_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_RANGE			1:1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR1_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_RANGE			2:2
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR2_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_RANGE			3:3
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR3_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_RANGE			4:4
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR4_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_RANGE			5:5
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR5_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_RANGE			6:6
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR6_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_RANGE			7:7
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR7_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_RANGE			8:8
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR8_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_RANGE			9:9
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR9_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_RANGE			10:10
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR10_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_RANGE			11:11
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR11_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_RANGE			12:12
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR12_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_RANGE			13:13
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR13_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_RANGE			14:14
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR14_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_RANGE			15:15
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR15_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_RANGE			16:16
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR16_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_RANGE			17:17
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR17_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_RANGE			18:18
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR18_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_RANGE			19:19
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR19_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_RANGE			20:20
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR20_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_RANGE			21:21
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR21_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_RANGE			22:22
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR22_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_RANGE			23:23
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR23_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_RANGE			24:24
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR24_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_RANGE			25:25
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR25_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_RANGE			26:26
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR26_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_RANGE			27:27
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR27_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_RANGE			28:28
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR28_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_RANGE			29:29
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR29_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_RANGE			30:30
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR30_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_RANGE			31:31
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_SIZE				1
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE0_COUNTER_RELOAD_0_ERR31_RELOAD			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0					32'he060
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR32_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR33_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR34_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR35_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR36_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR37_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR38_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR39_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR40_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR41_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR42_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR43_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR44_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR45_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR46_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR47_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR48_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR49_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR50_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR51_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR52_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR53_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR54_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR55_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR56_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR57_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR58_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR59_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR60_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR61_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR62_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ENABLE_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0					32'he064
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR32_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR33_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR34_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR35_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR36_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR37_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR38_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR39_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR40_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR41_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR42_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR43_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR44_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR45_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR46_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR47_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR48_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR49_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR50_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR51_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR52_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR53_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR54_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR55_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR56_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR57_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR58_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR59_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR60_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR61_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR62_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_FORCE_0_ERR63_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0					32'he068
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_STATUS_0_ERR63_SIZE				1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0					32'he06c
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR32_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR33_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR34_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR35_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR36_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR37_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR38_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR39_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR40_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR41_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR42_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR43_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR44_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR45_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR46_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR47_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR48_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR49_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR50_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR51_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR52_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR53_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR54_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR55_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR56_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR57_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR58_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR59_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR60_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR61_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR62_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_INJECT_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0					32'he070
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR32_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR33_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR34_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR35_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR36_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR37_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR38_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR39_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR40_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR41_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR42_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR43_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR44_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR45_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR46_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR47_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR48_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR49_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR50_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR51_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR52_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR53_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR54_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR55_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR56_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR57_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR58_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR59_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR60_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR61_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR62_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_ENABLE_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0					32'he074
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR32_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR33_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR34_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR35_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR36_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR37_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR38_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR39_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR40_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR41_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR42_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR43_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR44_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR45_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR46_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR47_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR48_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR49_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR50_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR51_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR52_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR53_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR54_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR55_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR56_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR57_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR58_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR59_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR60_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR61_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR62_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_FORCE_0_ERR63_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0					32'he078
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_LATENTERR_STATUS_0_ERR63_SIZE				1


// Register NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0					32'he080
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_RANGE			0:0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR32_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_RANGE			1:1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR33_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_RANGE			2:2
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR34_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_RANGE			3:3
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR35_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_RANGE			4:4
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR36_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_RANGE			5:5
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR37_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_RANGE			6:6
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR38_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_RANGE			7:7
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR39_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_RANGE			8:8
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR40_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_RANGE			9:9
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR41_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_RANGE			10:10
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR42_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_RANGE			11:11
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR43_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_RANGE			12:12
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR44_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_RANGE			13:13
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR45_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_RANGE			14:14
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR46_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_RANGE			15:15
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR47_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_RANGE			16:16
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR48_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_RANGE			17:17
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR49_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_RANGE			18:18
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR50_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_RANGE			19:19
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR51_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_RANGE			20:20
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR52_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_RANGE			21:21
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR53_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_RANGE			22:22
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR54_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_RANGE			23:23
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR55_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_RANGE			24:24
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR56_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_RANGE			25:25
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR57_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_RANGE			26:26
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR58_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_RANGE			27:27
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR59_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_RANGE			28:28
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR60_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_RANGE			29:29
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR61_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_RANGE			30:30
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR62_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE1_COUNTER_RELOAD_0_ERR63_RELOAD			1'h1


// Register NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0					32'he084
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_RANGE			31:31
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_SIZE				1
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE1_MISSIONERR_ECC_CORRECTION_DIS_0_ERR63_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0					32'he090
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR64_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR65_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR66_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_ENABLE_0_ERR67_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0					32'he094
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR64_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR65_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR66_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_FORCE_0_ERR67_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0					32'he098
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_STATUS_0_ERR67_SIZE				1


// Register NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0					32'he09c
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR64_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_MISSIONERR_INJECT_0_ERR65_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0					32'he0a0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR64_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR65_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR66_ENABLE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_DISABLE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_ENABLE_0_ERR67_ENABLE			1'h1


// Register NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0					32'he0a4
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR64_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR65_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR66_FORCE			1'h1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_NOFORCE			1'h0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_FORCE_0_ERR67_FORCE			1'h1


// Register NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0					32'he0a8
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_LATENTERR_STATUS_0_ERR67_SIZE				1


// Register NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0					32'he0b0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_RANGE			0:0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR64_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_RANGE			1:1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR65_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_RANGE			2:2
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR66_RELOAD			1'h1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_RANGE			3:3
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_SIZE				1
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_NORELOAD			1'h0
#define NVDLA_GEC_ERRSLICE2_COUNTER_RELOAD_0_ERR67_RELOAD			1'h1



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_GEC	32'he000
