`ifndef MY_GLOBAL_DEFINE_VH
`define MY_GLOBAL_DEFINE_VH

`define  DISABLE_TESTPOINTS 1
`define  RAM_INTERFACE 1
`define  SYNTHESIS 1
`define FPGA 1
`define FIFOGEN_MASTER_CLK_GATING_DISABLED 1
`define RAM_DISABLE_POWER_GATING_FPGA 1
`define VLIB_BYPASS_POWER_CG 1
`define NV_FPGA_FIFOGEN 1 
`endif //MY_GLOBAL_DEFINE_VH

