`ifndef __CSR_DEFINITION_VH
`define __CSR_DEFINITION_VH

`include "precision_def.vh"

// csr
`define CSR_SIZE 1024

// weight 


// input fifo address


`endif