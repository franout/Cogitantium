`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZeWaI1V646o3lfZMjPhfRiqH8yrcBHqB4Jp7GgWhFHtbq2FZEb45lF2y+4Z7Bo3p/Fon7Fuwxi+G
pfvZm/J78Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U278GGzuHpvR71v2lk6OfCq3UHPLemHH7G5nzQnoPxdKrkBUaO2E2nmWqUhjw/5RQf4sL7AgK0YU
DTyR1Zy31V08/arF1j8tyQmnhukfOHqr8ZKmmlkjtKowN6K59DPDDYpttGbqfNTx6uO7nzk6l1lS
Rsl6q24TQbBd1uaLrws=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pi7LeG6/F+tmgR2mSEDwUOPg9J3vRSMXNe0HxNeRq8mOvIHmaT6ypbEm7FgHQuSGN5PoQE3fMyP5
X1YruG3K+v9yk+bGce8/ZGbvghS7lU1h4isgDJ3niH+ALesIsr+TgonGh0Ol+XSo12YtX94alzmU
tkyr2R4bVkkpBHvg01MOuYc7cUQmHMBcy0p73aiGohZR42Sd4JJE4Dpnes8bCg9WMANMmBRrKs71
iPhWfZ8+p+ZM8j87IIQBV3IkpuHOArxJWcVZ6gR2w03ClBv6IOrJWD/WF8NZt0cfVRUoDc2P1DKB
ipFw8lJbMCDmw0VV517a0HsUZBxeyn0muuNqAA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bbIwBeNnHf2J5T3ZQluXrXgPlj6m4gdwenpJz3huRnilAqUbGa1gu2UEyWxzy2E3PV89zzGxuQ4X
5cvz29rO4f7FEbO07WMfFUcpIbFvYSPlSxQYuI7XvOEQ9QYMYsv5GaPrTyG09kYnpcmfHVScrGq4
pn30wsMt3ZIgV3s27Use9okvsfsLsQIc5o/DZfpI1ylOLXmgQEMl8FjUBSUNK0n4n7Ejtg4spgqf
a2jc9hq8hDzC7ukBc+mK0rNoXxALIE8Vm25bBWNVfkuOFKYtQFBlk40sbLvePUn/8g5ycOo4+tvj
nxb/oaG7tMKbswgJQIf9YUQoBcX3nQbsQPYmNg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h2TYH1lUjXbalHf8TK5hkjlQ30ZvEXKbnsTIUDUriXGbkyZM7BifousSvZesivmr3O0Li1KtytUe
X8B6e5QJLh288DLxi2Feje/jBR9xUdfb7uRl0Zqc/mkhMhc6PlTYP8kRpJlFPVYiyLOb5/mR9bKC
hI8t1lTdQmI8JQS+ncVrVb2xNCZ/nSnUK+AOD+nS8AFXCCJ8fs7X4HdDlmZnjcvSJNzc2pceLJ7x
8ADHhzA7/Csf6km2ypCu6k1ULmaRXaMQJXIpn1haQW+TNmCz/vj0i4/KoiStAn8OMidEPBEyG4CA
KCJ7cbm42dK7pSPjFEJ2zxPizwmR86ozsi1aAQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QlIHhNRjpFN4gXrZLn4iWrP6DODrKGhkK8sIm8VdwlCCNZhI6sNcceCfypEpeR1jiHjUiA5WpTiI
j4iJiEYtjpCbETgn9WkO3nceO2LgCE3RyuOgDABhkrAvDiNFeNUzgKquAEgEOo19rmp5ea/jLvYf
vE2VK8ql8jfwPNBfh90=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GF6UgWS1K/8tgAYNZd7orM2VWyBHqwif3OcunBF4fsKaVq8/BzcJgW0FVVikxOFOEP9MXjduR2kU
ECsJ8vPQoVz118Q5BfR27i/hgHlUKqw8/t2t9CZLbTAokB95982h3WFvO4mhHfqTwne/mCGbOVCF
VULMF7F3+LpRfYHMeplTyu6wSV+Tocz0+ohE9L2wTxo28h77pdziM4ECJnzlK0fdV02EbPj5Y3Cq
rAJHz3xHysVTuB5OFgs74lCJ10XKGk9d4jXBCMT9BJu03xDIgdbml/2DDg33uFpPPEWvO4ox+xim
HSGSORi0muLp9RWOGFqi6FFl6nW7A2EPETDA+g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KCmYBToXpkjbWHaI5FWDbAXmGo+FM7e0dkhJ+0ARnR9H6w2VEVRm4XH/krsJ7Z0ReGvxHW+eYCz4
fV+TxB5V0xo/1ByEcAJCqDietScNUOXBdb1CvV2rS/kgV3wF7gh806t8Dc1GLpw0uCax4AvMI/Ai
KbGWKs0b6XrAU9/d7z/MahC8ZFEDS3fr+P87oy1Z9dRlKEb1TzaGE1XcxtVoRbZ3e/4v9lnz82TY
r/f3iSMoRNf7X1S1UJWJJjOoMWxojPIesZ3Y6lYMgw5j+wBIfS4M19hlYakoPRXHEiJZVvyra2or
G/OIjuk6GNexumwfk+2MOEZ5ZooKFMxgjRxUbw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296400)
`protect data_block
VxHWHvmmw5rttDFOS26DXNV5iXR7VxbZiFLx8WNu5eMoa7rJgLfhivDI/WZT0z0CdB002o2oQQxj
ya4fOX+gz4DT8YwRX5HdJCPrqWH9eNMDcb8U05+dF5qd11D3w1qtldcHuXNYoZU0wFlvrOSy04ZR
rdrwrX7wBMlQ9KXtF6p+8CkWJiikKji33aO4MX6Z2uRxUwEG/tCEVQMNctEfS8Sz2s6LRILeCvhM
gscPjYOchjcXS/r+h+HMbBgOxlVDrArnPgViIcI9cdnVrrMw48LXf2BxgGgNaug+ZB2Zt9qEiOtM
zbHbNfSkSsgAF6FlQX6JaxkaelEBl/zl45zBH4rAytLtyjCq84Qb6q6D2iEESnqYRzKh017r2QLL
/hJWXaJ+ewobpWKX5CBaLHFsWQmDV3RakHBnAFPu0zZvO8VnG3OKfDfdVTBxle+1rTwQbypdvHg0
34/zXSt74KtDe+91KSsYpiLXqVkwDG+56o9YAdXoNdv7f+PvgPfH02UbjIKTHl7t3eRMg2eiv0cc
ChxZbBpTxXzaNPg0B6l2Vi42/TsMX4Ec6iVaGE4e/C1Sb9SYT4byev6uPHbrU0YUPIVK/2wSn0HQ
YK6BLhnfyFwaHEBqN/41b4C362B8fBHAZQ4COSNABBypPZpRK8PKGuVG6dGpVM7FInqgl/SN0MsD
Tf9Sh5ujEwy50gGF6qwBSiBCt+w/9hDeUSGG5w0gmv67TR4KvO9FxVCjkzDryZ+cVPbIvxFu8o7S
Ovb5pWVNUe1tm4DchN2YWYaDD4T0hsfmG3mpzIdlzvMK5eb/Ufnrfwfz0Y2VZDYnj4avAZV9hTgw
UWhDi/x/9y3NPK/cuZLEnivoZjPZvDx1nMKWMtTUcPCQL4cu5v4iPU/YghG9Uypqjv5wvO75OBH4
vB6Sf4jeAhhQp6N2XI0L/5XKxPrMfvHe061xv664C69gVlRX3hK6sl9p+dQP5jOnZgo5/04OeFcm
9CjUPXrw3r+d5DhiX0tFPwEJIwzCWswAcP+eoWG0WeWzKUT2QswP68NU6RMWP/H2JWtGuw3N2Owk
Uawr3inRxPCpjipOza0aMX9Ti2csIKObMfdYqX+8VcaMaqXNpd+yFPa7Nph61+5To36lTliUlZ7m
HPTTrkDU8DYUS1xaN4Teg/QIEAQ7O2LHAXdedJbRbedWOj1TX+4pdlj1YyJt1V0nd08UTAXBhjn5
FveBbpGr/5P6WVKPQbQ4GobVsNtkoQINes2sHdWSLkU+wox6ahlMboHiqxulMmrMikmy2MgkAyId
tayK6jnYEbogS2WsTy3o4s4CxbP/TzEVfQXtCUESI5r4Ifm6UQ8NsPiIxP9McBx+Tt8eNjp+f41J
IHruGzkTS5hisXSJaGm8mTIyS82IJLvgOvs+/O0PiKKWsM1DfJwMrPTwBlBtzANEoGoAjXgD/D3R
j5PSKI2znbM9g+N3cw/q9JzfrE75exxxCguKpa+52Be08PtlKFpQWY0ByUCXsbgDUiT1BcXT6Ocw
15zuJRXhOjK2A5XGLN/TigWBs8urA46O4B+Lx8+0gvBABWhb+NiedtvEsHvX6baB9KKsJRbJBpwL
yHufWLK9/7eeipolFD2qiZ4q652RWEdvF9p4asPVIaJC5QK/qNJakbI5hx/pilTSF2nNTHXyAEBn
6PGVhviQO0OvyfdhoENNfnkkk+jQFx9OOfGqa5bkyrvoK4iuvjvlKvWDVF+Y5dFdYReIlYcn32eE
hfZyHRYp+V+v3NdpPCggEIqYTH1X8z0mVD6mPF80pGfp4qF664fOC5CaXGGXkwAHj4zREkPs4zg1
2OsYYEwG6HpZXd6Bf2d23jeSRtG8bU2xAulRNn31yq6+wzsaDSRAh2sON7QwmDuZLBezhJw3kxJv
O+5mQurGFKmpKm5j5tp9L4Ys3LG++58xqh9tjaYJSf7TDtLRcC8MUjLK62oQYVajX8ga0wJZ9nXm
fDR0kQpXBMfrHyzDihM23MVQ0a9OSjkXdoeTpsOggHfv05iu+r/RQvvsNVWVf+2rk9tgd6XcZ4qS
YBXGMjdtJjIA2mWOjvDWlYJ2xgswl5+Abu069w/CEyxpkXUZU9B7Ece3uN6FtT592yrwf5XGSs/A
26w6/SvM3gxS23JqfbxKePYQp3sHUh/PgobU0qOje6SGpD8wpKYPEsNiFiX/+7u+eDUuA/3OkOO4
2DgIdKMK1CcZkNHpg/NrCGhiagNOrydXp9SF6Z8/MvOb87vXDPAXt1JJxJC12P18hj/ttNabr6AS
IqIVqJ1X9nXSgCZpvdgvWF81cwOogQTOkfGPsTRqxIcoTEpDkwRw2399l2lJMIptgK70X8CEAzKS
1JX5B/2iuEyaTymdXrvdeT/oShmzF7t7T7DagfI3Ys5de5qDNIfj9/4IIL63Faq6Ukb1cpRtiF2S
0xmkE0IlFDC8huKOFmMabcYZaU8+VVJa6CTnckmPtSQfOkz3mzH8ZOToypKapYascXfCLAsvL2eE
7Ghf9UOfmn11CjLhG9wcKHMNO1faAqgbtis68kBY7RJxuaGC50Xdr0Z7su/+F9UfvIi/yAwiE4H/
nfze3iFfjZP7Iz3tmaF7sDUnutZjaCDEu4UxdX3EqUIFHB06EgxomneN0+lHWDU2iZlP0PYmJnqc
8jqUMeDtQyTnuXDhkFY5NSoOfAgKoiDUl1/x/tebAlFXq0ylSCwHGj5XHVb1uT5vIZM5a0lPk5dE
xwULaZUfWOmHo+wSXHCta0+agzluHZpMlx4t9Qkg8UUnIuPzXskkqumtOOnqpCh0tQUBQUOx2iRZ
PgvQZuU1zwa9gDOzAdmZvISCEfJlMe3WoM3dZk8/dTrpNs3RZlKD9TciNNXEIMyyhC9HdW+OOAmn
HnZ4esS+zqCEPV88LX4+keiZFjjVbH5pfyZ3QHgd9EzzNsufwHZ5WA5JU0EZv12Uipf1uwxthdq1
02PIXTtOyNjoFdmqk7nNZ6LAfvXOQy7wblv+YxBATALIMYkWOe5ZP+b6w8TTwFtV9V9zmlx8oPOy
dRCwK/WVIt18C7ZccrORkHANjW1yR9AMsnkS40UzCXXFN7WbsJCoFsEijHptUhnko/VqS+1S9YmB
P88Ijia5/8KW6Qlo0K4ghX8gNBWKqlorFS2SkMQgh6tVxh7vd9feTRZAhMAR1aW3omxYzBSrwdw8
1lDVW8f+LSfLEpHB+jMXK9sJ5uoDCsK3Byf1tBzn6CJ7eP0to1L7z2TwMdOlXshvwZ5ykyso8cNS
iUHzn7NXrOqHXZQcbUCRAO+OaA9TyzlsGFmsat9aZZJzCfTO/j2ucohNkA4QCxMA+XuMSzfUM/Me
UVuqEJUmGqZgcAhJMzQejSZJys7eeX8c7GcmkpS4+gc57gRCmwCe9zAWEV6n21Qtl9+Q4KIpd+7R
EnVN+DRrFXehrX86G1U81d2YYYl8DMzh+5b1X8hHsAoS2F+8Hkq5JGZ23lTKHoLkYwU8eXqoplpk
bYGrjoRQ7JU6UYDz50NkSYfggR7mm0FtZVQaHiqfEKgJUfToCUj48utcgiOVj8AO+ClsouI7H/O2
8jwG0TUs6kPXC6ak8d3IuC7H97BgWAaOaK++/LlfervxU0LtU6183xYlrDHpSzzk9uyPAbpsR7Qq
G1rbXQ/G/GdOsCIyBTlt+eKZS1XngyXGBoM/8Al4BfrWyEygGFXtrP8Tb2ZOx88V7hedcoAMcMJO
WRc3EOO5p9LlrRf4mXWDbl/NAI5iQZDqj4qQ9JhFRw6Is0sh5yGPBlOtmhF7aikKmondwITdpD9H
ubY/wLth/Cmtp3T9jz/09dBfFrBcwFUgqvbDBwpEAKfijNdhCUxCIaIVVpBnePVRUzpqXyOfLGfq
ux9SRcOZ/UUB7bVudp3UZqGKcBkmZ/7u3Mi/DUtqx8CuNmYEfNQJBB4bPG+z+lPWS8+y0e6FgU7E
YuWVOLaxhOsBZhqpfm7PyENeFIlFIfk4rN3irLpQdaymBnlxMa1o/6N4JIHr0C+cqD11CRu9i2t4
CKLwZx/zXXWY3Ad39eD3C+wSDSJFAU1pTcsbW7H+s/iEYXsd3hZcOrBMZj5NEcjvDHxgvORiOevU
PxmR5zz7Lw4NQfMqaVfJ5RuvBrNNtva71mjHGptFBSR84zwyXUi9S1fnxo1XT/1b38hk5GSzC10v
NZ6LYNr1HsgbenLxt9ZdVIwnyZ1HdgurOFjkW6ljFcVGRGZK5OJYT678bSED2eo+Dn0G7Yij5HW3
+iQUHDTUgy4uNSYpmlmFBlKtg63EdoSkxs5K/oXV+llZXbWodrwz5mIqixoDBwAHaekmijBAOKci
rJmYhK00eUJtH5hGfPEFhKwTJooSSmjMT17rWGXjJVXG2Hi7YWyj5IoEjmohlMx6yJzxYhEPEFIe
YUTwGeZZjSgtnf4f1OyVmYq46lbUy+edcJiiM3hoG6dhuxAujOosAkIQKyDiO9mT3d+LNIuO5iR2
RQqfFaSlsdv0B6afxjLVcX5vLRF6QgSGJuW9qBJCV1XuEZSZeb4LqNpWaC4WR1Kjo9odXsSPerrg
yriJpZpCs1wlbyPUbUjKbMT7BxhH1WnU+/iQQZdks9nncbORM1gBufJ7T9gMijOldEsMfEKyhB9y
sc0hKvmH7sdfvB17VPVBIQAmFfPUXVhlrRJK14LCOtdnT9Hfcfj4EqqDB2YvZNV26HUK0DIt1sXS
3SJEtmoEjfJbe8k5l+mhYTTFkr4D5vIiGOXf+0wP7j5NbXqoD2V3P0ZP/ISLtoKiM+RkXQPYt1/A
kRNPP0Nb1v09etTNec6Fz2PzmHkhltkAIls8U6cDH9g/tBjHUvqrvIMv/RH6KkwUE6SIkcoCrOT4
Z0UIO6joewMV0HQAT8OXuGjNdQomrsvu6QroXzk2ve7E0p1n9mAv6te3UJvd8CCc0MSsmrDbll67
xjPv49XDiarBrHtPCzVMLk0bSsig9t6Y+IYqBAOYhqEnN5l6GhCtZQiOtO9Yuzs3YZOi39ji2ca9
RFurAvuY9iib963f6IF/cOF5VtTyJaNS4tuhLFoVuLi1sRQ+7behgOi+7xfPf6CZI/MnbuJxxV0H
gA686DOQHVeUGkvygjaKpDL0he3C2NeYOFmQJVlCOT8JzoFj5rJ8TXED00giFoEm6AuLr7b00xUr
bNHP+NB1A2lgcbsbHQBhyVmvxP+4fPEgR2ZrjnAprW5gOPQEpy6ktjLJMywfjCG0ommtaUKM8ab3
Wsaw5471vyTEzAGOgtwSGQ9RaCIVbHa0ArrZ9x5Z9K84gpVINw86abhZfG0zp48ysgmOWFSh6F9t
vyTpft4YDb4VV8deIinCOZbdBUBDtEtDb4IRkv1JGlQk4gPmbwghi1HMTex+H68SoDrqB98IVOwl
tw1iejCWJufzHAuvS2KHT8ysFfDu7WI7y0znugKE++8420wcZZexOEBpzqsFaWLQbMIrCOoc0D9J
dU+tPJh7xna4eJ8WmXdNWpZDzFRCoT4awH3oeUOBpnJjk3eML6uStROrBdQ8CAEwvQWFPgnK0aY1
WJJhyDITaWfaoL4lQ5xGeBqfyk66TtjKrm2sIxkhlFHgyZN5TuVztGv2ZgYqIV7IgxhCPH/0ZtZe
4TBb6RYSmazsg4ufyEb898fpyPNN76BI8rh6KjpWWiMWGldJ2SFhWmCJyb7bSF9y5kE+LAv83DfA
FphycbcvQSkVexkWY+H7tb5/DT3I4mqmVZfZdGwNbuCNvP5x7NrC4Zo92dWGVWWDzGbDuO9ybBJY
LDPrZPMsMCZ1bcFjXu+7zoeV0fnFalT8Y/Z8yONQPr4cxbUndCRcvh1A2fPPpVDuerllX/mZ1p4a
LVcm29zvin6pIxalNZLJPZp+TxuiCc1QgcBakNf1M4hI64a+qPZs689SpjCZgiLU2GT1VMlBp0yk
YV9D2PyGNo4M3x3hqYAirEwI8ITUnRC1YDQ0rMdObB90ezoDI2wy/3BAsss2nOsoq1iVgogIxjF8
1Ew2bCdpH01wByatKuv1ljoLmXvfTYpgkJl/Wn/viM5VfMOkDut47wnyeR02fQGGhWhXyBkm3wjE
mebqMlk/bSln9TdDDBfuT+oJvV12ib5cL7NEL8abwQH7hct6Ei9LSw8b/1/jL15FBp+LFIwfEsai
Gg7ofmzdrQjkhjBcZ0FlYF0l7F3nLYBjG0QsQ9RLiyGNQovJ85JR5RvJ4W4t/8Ez3wuXsxX4xQ4E
XWXNN2LEeVyleimQCuFvGggulKkc72qD6PmWblLvtl8VjT4sjmjb2j2mPx/xmz+Ee4/QywLEdZFi
inxRLISz6Zmy+Gj40HRx8q1XRh4BTARxWdPAHNl9KI1toOCTf7tMdpnk3IenVGVQO/0wo+ODbuwg
CPe8Vkb0WPEDSWiT9OOlQHWlwTVSkfLhh3mFVCHjviFZ5S/HZCJrcyJ5OZIoamqkr+2fbLPGpuNP
+uU1uqPweogbByR/3Vt5uGPplnxBK2vLADPz4iUVTIrgV5GN/Nl2KtMU3lbkYiuTf6PVz126tfIP
jOnihJdcirEUVqq5HbS4/7c84Q2rNC9zITFoX0QVR3R+mdCRFZC7u4FgeyaUxYsWErbZ06mc8Sse
KQw18TmnwPuGxQiMkPEmiOrT8ENU0ENgmkq+OMzPHh8CHKiWW4agmH30E8uApY8PA0VVodxco1lh
n2yHVVE2IQU5XfpjGXFgHjaz4D4nQJ1pFwZrZo5nL+VrRsux9JKBBRUbzMYV1/GV1VKIjtqOFqns
T9KpcH8wKVvcGTb3nth2yqOVRlKsJeM2+Oxr0zPFCnL8SwvyQrXYyX9+JMeMw/w1L1x3Hq+Psk2I
1B7jEmudkenecKAB62BCiB3W/yz47xa2q/u67vZfJIKasQp9/sarf30/Ucq6T2vjP+4duXqeQU+S
rfxICURmVmlZpYTBF6jzgmAQSLnzvHCG3DyZE7JRJL59YBAnHBWAlxA5iZ3OGscS4nLt9l0BlPAo
/pHuQmx+MBGL0vqz8oIenQCTA31DDdSryFwT7Nkh/pEaqEMFvJmeSFzUUChkNPdGI1ItB6gf+9dt
wIqZ8Tce2WGGQrv9GPux8Y/8PKBIiW6DkBstYiZQ0X6ZdpQj+JaGT0m+zBiS8c4P++LvIGDVgTJI
qSoGIX7J8mNUAumhNXDH+y8O7+TyFdDMwSxQSBx0r0b7La+X3REQXSPZ0wzAlLTH0OiunMgPuV7h
4yeb2oNikr1QVwiHLhZSMaWf0+TXTRDj1jSQuLlY0Xui0Vbtpwh/5wp4OcG/oEs27pN5EG23nmyL
+ZjnCQ5coK2cja7Fw4SXaxZGQk+7n7Y+jx+JDIcJLouObR8pv1B85VdNOsfIuigX2eEtJT1kJe5K
sUJQZOXaLybm2gOLgd0GltdX3GtTJIoHH0RYDxUUalWpKFO9jqcFlXKt2wADMGCBV8KTlee8mCkl
oysCiPq44xkOqL9E8GefHwSZkVtnZsH63E43y/8IgpnCGrZKJ4m5eFXuYi4HQ3gAFqNWpsdbeo25
XKkca7cAKqNZQU8nnBmkXwYOU+P5AoPjZxX3AocbeiJwe9iKNdfdTmFpjMb58F5S4ld4a9NrEVux
0Bz2jFXv1D3U6FgsQ0oZyY+0x2fHlK3xzowf/9LpuI8emziZKy/ndR6BlP8sKCUNjt5/SbKaOEAN
/oeuM69due4TxO1tJFtDOP6OzddDlK4QeesUGp6UDVcEDM/maY7uYDkwht408WmTFAgdJas7bML6
Nj3aGLRoUUZcWF69vZAJOXUZpb4cMPibCEbRH1vqfBD5d32HHgALNzQlYCKi1OxzaeKbN50ElHtk
k6/wsJWXkFMkFJAVSiDGP/H98GZjSZbzGwBPrZmB084BqEXBgYuPJ3VwJkWFqGgkIJb+YZNzUAlm
Mp+59lwCn97vJ5EocYFu1q1CXGYqkjHgekjpEYU7KWR0AZPK+gSNmPNSzdFEaGOI4esbnklrIEcb
bEtondO8rqbA+twvB6SOKK3G34rW0U6lZTLxAoPExD+YxJ0BkTMFCuisJeE3UDTQBBDCRVBVqGw+
SXvrNRu9pxSaWbO6jj1b/1Ps+FUhzAlSeUAGOvKlSGS2b1U2piuhg2qqVpEiGVRuOgk+uSoDPtt7
/aKSep+6jmXpYB/aRxFg8/NWSbEnvdfeCdkFT/0O5VREL9IYjaq+g30/ru3j44HKGLoomU9Joqx3
wKx/0o6GOHc+EiTy71+iMad5U1y4oM/jgj0apBKU8xBFqObmd/W0YchmBX5ic0qeosciI5+zjYxG
VzMxKxJN7cMN9hfcoBFTp6ZVBJ4WXdycXZW/s+lPVyJYiZXhCH2IsJgkuDhpQqiCYGPUMTVw8jx3
ZaL8aLjqn/xx1BxXlYaqe4H6jkqMW21UYWswWhFk4W/y2RXu82pMeqZdbTHIiV4zGucS5H9VTg9m
3FDIVBQM4YxTvQWybIB8DOzTchVElqIzhSm4Y9TYX+YHuMWs0aLmku/wZ8CtY8gRAG93hylaqNQ2
u2fgbXaKGdLT6YQxL5+97BypQik5Lu3p0jf37KO+evRcqjzeSO9sKKWGdXQZyBa3R09habwKp7+A
io9oSmjqy8yzY2+VOY92rKuxGtNPbKAGKpOelRtQJM/mQy2fybB3nU28pqk4J6bgQYbC4awVtJKR
Lwgj+HVXc4C5/zYMUsQ1m6P9c/wH2gNQWpk33rBToU98gnRbRki060eDOKGCHjvQLwZFbGhXuHTC
6IYzIWvxxhRVGU0011Lrn3N6BtoqJD8tk6Bm5aBztDFsBKXJf699D4EbiUtH2LE1eFCIomNzthVi
bINogbK7U+w8dnzlLIO/GaMI0io18k3uQyW+AOefNqSgUC6x6hSiTRkBHYN8EgRKZjM3pJ4tGRWE
kjWFCEOQsbOOChyR58y9io/osCNMcMJ/xHOwTQ+7VQAixr1T3ziGaKzuD5yNtv18gtUABmXNkgz0
DXCqHu2IKbA/LdYMN8GkYJ8ViUxiuyUy8+U2AowPUdLFMI6r45UN/VJnXgds9IEHupU8GdhOJAl7
SvKWaYPfDhjXLbMFRBoeo55cmaWIAceZXUgrE+H1zB/jEN7tyFJ1FL4W8xO1qrEoUOMgK6Mnqf6X
1eVYzirMOuOJCTLD71ypsRpjyJZJCkWSb7QZwlqA/Rphsdqk0m/JzFovuLVxQob9+XQiyCBleLvI
an5vBAcKCMIjwn235uE7/YhPiMO103tGUKL3Rk4J/d7A03UZAbzCkTjviVVCUiixrwgTAx+k0eF1
K2qXbz0BuYEhZAoGvwfQ9HNADbsrXrOABji8FknW0Mcz8REka2k3whesCa8rrFv/dgSzMxkexmNJ
g1Ijnn37Ck3VVo4X4R3XXZ43vc/D5R17qI051V6ygphTuo/E/cfD/n7gqRm+rNkqfvdaWeeqceoS
DC/7grxEHUGYy+uTxGn/paOw9wYQMuNoCxKNG+N9bXBjYm/yOJ9Q73227ypr87XhbAuRUXwD7ZyB
FhJsxoz9Ti5L8pB58WH9w97rt7i0bHUt0P6iJNNHtVIhqHG8c74A1E7R3We1sFt9thPTRyDz/qNz
7+URS5Hk7nFFnxQssEF7pbwbaHF2/QtM9s3owXVySDFvQRSUJiQwiKndeWXhGOm4jaDsgJJZcM9u
UnB2LAdYHiucens9GJInu9A2kc1+ln8TQ36iTSncXeYwvlhGYgRwpF7jwuEP1WVyuX6uc7nMPFCL
FPiVskQBmTjLuGKJ8naQIl1ErJA+AWmEbWdq6EqKnuMb/iBScEL2slTby7y1BKNu+cCQPmK4yFHf
PYZ1kex4FwdLbbiFGTg1Q7pCLT/fhib7jYeIv6LNqyG19DlMem4uXsLAcIRyuI1AwqTB3hc3nDAc
46/eS9ipyw1r/GFsvAVsFh3+ad3sbU7ZJ6OOHbLaM/6n5kHHOt8/Inagcl6yLJ95ql9IAwls+s2V
uJLruUAldYLIrrIknQ9L9/jYZ6QUYTk25AfVaTgJa2R1SVtjfg3ALlBGZEyQYTeTp9xctPGzeXPH
DgiLy4/m4Oepfe9PlxoSyE5fLSZw/pRw2XO3PT5Y18nVCF6kBrWRZwp9Io8ujIrkwjM1OVVa05+5
sSfkVjS3nDcPaC8jZW9lT+YANqMiW5wTbrvX7yrF2zsVFo5gpGqKtvK3cw3i+FHAbmL5bUYPSySB
68btXOy+dpLitwt+FuBzGL5Pr7vS//bJ/XdxzjPz0S8zU4EcLajdMKVh7+mzIUw+7JMI6DPYuGIg
sr4nLuBIFyW7YQJLiFPvM700EL7Jfcm0Lht0DyG0mRH6FQ5Qv7gegAGnUPcuXKRIjlNXQsnt6Wd3
NAf9tiBCRGyEuE3iBj51UhAMHEL+uJIYLg6yAAJlSg+1Rr1urNeM0L2ekNFUfAUwkOnthiNeagp6
yUIeHms5K7d3vIb5YNu+c71LgPOBozDg4zHoNaSoVA7EkQ6fhrpEEhe00yhQqppiptVlw7fR5ugr
zEEFQg8DPadBp2/nKGo0pSmqWN3eg9th/rGoPBcf3QiWszzRL8Oogyu7CBABwgYQeDevfMYD5n3f
pHIGpZzaqNUJLHQECfjGwZAw94xoMw8TbtQIjNnr0hC1GJ2GnJnveSlVvCzygLxFI6OGJm9yM6rG
XVfjW2tumCEM+1A/ZcRF+S680PgIcsN/MdexBjTH2JY4rEY/aXt6h+4BizbeqqierF6CezTh1NoF
JHODLomtdMH/CK2zolM9lLnlv0DbQPbm/OjERxogv6VIFS3O4iqQ60XXlcuT+W5VD29BqmFsGuFi
u5rSbLzc+l6r+VJ2P+61hpBjXP2K7OiuNoDHCO2Vl+oMvZlKHCuNk76n3CWNQZOWvh3y/oJDIcTd
5Lv+mCWDtfIQnCwWpodNuUKMvlZtWi4Q3AaDxCo3EhSb9pB+j4OpECzFIYVXbUB/RoXN0kXnqgpp
/7RjOLque1cKbGE1pUXO2YPg9v0peLCGU8pqC2YdiIepwtycXTQKd7GA0TC2C6TgXPgWXodtdLrb
uuV4KF2p9/UbTxQ3ROPHYoLzp/9BZjiyQrZyRvkWLlNG5nRcAqX/ZTc8G0kcqjNJ9jA2IiJcT9/M
pvDY69EAzbbt0CmWWQARNKPirq9hErQCisKicXBpoVY7UdMDYgXYTB85RKEL0TaHaxJ65Odw1q8V
bE0S/knU65yvSOb+jfhmzhvKkLSiFXUdOEwA9rnJLhd2HCOzPfAY8I8N3y+OHHE0Y+4EP60tbOxN
Ad0yDuoFy2k337H5D6j6mQXypzIJQnjFH60wzSB1kawHapIZNBW4+gDJJDHh1FUkTL2zXzEI7Ckd
wYU37GsjMWSOB16JfQQ00tM/0v99tTAVlmGWldChEUldGtAIy6SSe8neRQ8QYVRTzMC9i6t60yJS
ysbz2hQoUnZwI1GDSWMPtg4h1UDAk+FtY0IoT6/4LHtBy8s/cFbgiT4mVxKXxvJZbBuUECNvrEw9
6N1joL6m1XeP11a+QXKhOgPVeIgvARm2DfLZYhzYAirV6Wy48YzspEX+UFG3/0KnaY/kZg28DM0i
P4YxYYNZXwkw9esdA3K9A/4Jd5vLH8OAdsWLZgEYzPPtG5Y7F+JOAyadZ99v8jrzB/Qbd8qjTsjS
bC/c+Y+sb/0Wssi5APTvP2lZDXl7Au/7NCLow/IdTBmbnMNDQl2k53xLgqfRHAJGJVw9X4fX14j1
u3iqgUb6UtaW5EDLz8QHKYNFntPSS0F+8K3Mz8q3s56y25ZoXYjgbApdgKn7hrn0HGceczM7B7+F
FDkBVsb36iJKs8h19hcjw6MaertI+9tB/P9iUcmmuoJjedeg1DItgaBp23strKQ+CA0IFrvCz4RQ
IaU70USwf7xTcf1fwBJePZ9GqV/5m/W4eiyAJAfinzpL2g4AV/vbXwl1HO+lSjHh51TkQ92yFk9z
OFQ2i2WTc7RlYTlVl4ZcTp6rQOTTpQuW2uyIGTuBA09yfG30qlPlN3npW2sOepIxy3thKg1QTfao
kMSPR6x4UfWXR6jdmCH5lX73U4j8OjKWRdiUWYf8Vy8hSuK34e/dN7H6IFsyKLXk8EpUD28SfUAL
gd6uDEMJfePT5egmZgwVoX6jAxi2nMREyLKdaq0yrvt5BeUs1zBpConseAaXQrUfxvZPpK3OupT/
sfdX74ReN2tJzUaTPt/m9B9YtK/JPn3BlHcRJPqWu7LyDNAD9E1UmxIK5bBy1ajdaLidIRujEGAP
N8KYpLAL7bRE5YuKC3rzreuWvS6vmRrcC0XpOjk4Rn6x5345FZ8YjIkQM0NgF6GGStP0cvOTB8S2
NllevXLaQHwLD8D57S9y/rAKHAgF7sBm57sEwpwsAaIcVQamUewEByL2gf08OPzjIuewBsXdQNkr
HibMFNyk8V/vBw38YKMVKYnzdGqxEdOnvc9E5yx2KdaAJyVsbOwHo03bht2L/JF8onEtEiXD4+ff
tdG7f+ow7FR5UEPhCz0JvAHyEyt3EaERQVFfebUXCMlXiL7XniqFSHeJHdPSgA6tA2YYLL3fv/1/
WEBBBJrdzzn78uEUVSIN9XAUNYRNSGRG+AnYvIxQf4qBlfAs0DJnoRVx54ySuR/Qlc/T53jWBEFL
1Le8s2TTGZgnzzS4btgGAO13hqpfgPUnKyU4CQ9l4RyKXffDJj8gBKCYQuN7VjwNlweBEvhJrrOL
RFf2kydswihltKwqYmyJGbXG5I540B++TZEnznLLJuEKL8P8AeDpIYf8rR3bCDfhxVQu4iOIMvvn
/iNUQUEP2PNCPq4WYS7g4iKH8ec8iw5NAFkvQ5Drv79tilmjLE/+VRUi4v5Q3l4iK+rOZ0F0KR8g
oTFMwlyUKcLJbCffeI+C+BVobxfLSTChUwlbYWC/T0i5t7ndBwakpUOu5bahm20CL0OiyBSUDpge
qFOfRFsinBowdt4+q6gWrj89vpgS1vaHy0pityLoPxT4K01iRyzVGWwSlbSLo7xgeXzaNahXa224
wmlaOS5lRQRCQsfjPcSX41+7I0Lr2QzToqRAVJmUSo9hbUFrvZT/dMH+pqwNEMn/7BZ2O2f62G1E
lkCKftejdVaLHIkfNpNa2GdiMrGLWOUEnmS3tHBYcMj9KfMVIN4bmoqIPCZ3J6U8S1R2XAPktRvY
Qp/uz5Wg1H82wg5BLTFusRzZrnf8vHOCUcuFa1orPXAUxElAz25xpAm7eZx0qGNrlP5/S8K3SdYi
m2u5gr24dFPzeao6ymPAI9te94AK4hW/U/Poc/GV5Wuf7pXW3uBplyoej3TfqzcCV+0f0vwC7KC4
8HaVsoMoCkAbC//tkQFc3KkMz0esQ9rp2AFfyhIehVc0OxrYWmchWSxiMW8VgUaewHDgLs8XsU7L
mfRkzffxMeYNet1qy07dABCXix8m4Ank3MATA35RBhYknAoBol6exc1Z6MTHw72pNN1XILXiPyFV
DQGzqqWHqwQ6R7yDKeSJ/LII6VJadzMqEzX+6L52FfJ15F9i3vH+Kex6AZAsKh3lY4kfz8FMFBJg
BW8NOjRQ3ZnE7WZsXAzo1kP8g4YzVgXBQsBzVAaExGD7allJm2bxvZy3WHA/ZYWOfS1SrK+n7dHR
yXBfw9ETI/BcXF3VXH79mjKcab+ZAtE/LaXZltOKOvx+cPELJYQoHFMGCn4ts9Ba2LTYl91VLQAy
fxRI+BUra8Mv8OLwp6sh9XOZQa3FdDUmU36Hv0vA7ebre7+bR4Griu2KiMoIBFJdtqKfOqO4Ijx/
9sI8Ru8pZL58ZlQoabXAlUKryHasBQvtHmBsILsARJfFx1bsKxL24Qb/O/HfqktHNbeD6da+q+CH
oclV6QiBQTQk0jO8nTEWkHKBcWTsufJmK4cWMBMqGMqA4/tdX10rDowHBiwJB8CEEUlfFG6KAoEC
kqxkgDDT8Zovc8TlFMZk/XAA44qJrIdrQiuqgxZ2kC3mUkcdPKdOJSIvZVHv/G/XG+X4Mf9DHMKH
nTUn/gAn3sNmcSFjB9ftLGKr+IpDqMO9fdHy1nppxUMtTr8m03LhbtU0p70KtAvNQLdCHNF+ZJBg
C+myQVgSRTeflZLjFVg9L4TvQ4hRUsnaI/x8jTxgFg9pG2Q6amoJXQhqw9/omo5SW6h8YGKU5mqW
pEmGKVjd/R8xPsPxX5Nfezv9a6hC8ItIIpJmhhSgYiw+EOlhl4pO5wz0JK06+P6StJSR1M2NoqL7
rBE4nBtMzjhTH5+9qxsXm0q+/QC2rS1nj45lLJqs906UmSwonIkNAYVBxbbBBTman8PU3Hspm/Rj
p4fnQcy8vmoLiY8op3EXNx/EE37zw9xDzWLEm5BYRuIHaughFdCLVK73TZ6NcZfrdqSiGLxu/alV
APfqSxxqn3dGKMR3EBhA+Mdbkvts++aJt+6dXWP8AYhpBfi3AGVsibFn6zcH69UMvuEFMEUCLzAZ
61MGzIz7FdR2v+HBCFSoeP1Mp6at58/g3EHkQbyAnBnp5WbOJoi0qmRABWpDDmWigGRV3xk8oLoi
o9Zgn9HWIbLR2lX7SxXaBMHG6h/c2tqKGnHjLeov3ONIm6jPL50tNztx2Gs8W6D9AgTC993dfF8H
oEE2fR5MDE4cBNMrobb89zU60BbTpIZl8bfkuhje80ZbKJuHc61BfvVvINxDsOVKtT6hhptWBbgV
CQAFOtjv0gIpFCVUa55lRIhjbVHMHqkmHZuD7JpiwQcnvrncwhKHjdr3OKSMZ6EOGh8I7Hfgpyfe
/NOhRCRokfYBL0Kx8GNgaZ0W6q85njnnuZnRU9A/zXO0mzzJxYj1Zg/md5UDmZN6HhIv9oINwJCI
YWraRgXw+UaVTJe+1j3vTrJuvYV1XBYFgTqiWq6tDAn+OPSRgGZH/FbHmkaljueUImoc87kU61s1
2w9k23FB0hBTm3edUutfbPeoaccmWR9+pgy4WQpjxh4Gs4D5NdjgnA1W2BU05xioKFgJD4qJ2HqW
p9kXV7SfgaPcMNnx+ZkZuNv9tzcrJhmgkJey6cOzzgeebnFg+YgHKgLG63pbSk+kwh61mnAdCDBf
+qtRz6NSyNJqv0GxNx851Zj6Ducszz4VJktlEsh0Jxm94PxD4iPLRsWt6/fUE7fuG+sa+D4Z8pnY
x15L97NVpQ2EFR1Ujg39w5qaQVWbpo9hfbbyFE1RzODK4NZB6ZKLvjxecmNDDwywZd/sDb49I9nN
O/ih1Bd1ECVID1ON8wz6kKnPOphBIedtYDewFSUDbiRTFXAJ2kESmMTuglz1VDEPkxAYcVtCAWUt
8+ObTTI8LN+ojH/FR9WDKtsnltAlAG+vajSv6vi80k6YG9n2xaN75+/9bGn0SCIVOugooeTAdnj5
+g+BDeA/Ey3RhgduUIkF/wDIAhwMVw/yg37ePLUZeW6PlfpntIk2ifFo+rc6q67KZcNKjuwWaBET
B5916fWFzGypDxaAapxHoSHknM8EYNZfWUm4FmJHEjj3JduyYoIss/aIK5shwWco2Nk86KhAMsB5
SbbmMdcRhVImtT5+GxtLOoGGTuKFbe5yslpJW+9gXTDabEoV4kj4IjYKGuA4ywjsHryx5AzUKjSl
Bp1FI837kJ4+3eR9Jc0B4asAGHltO8h5FOc+9UvwjtBtXeLCVGzXgFXGHUUkNKlJ9BtWDF7/aA9D
PWX+3gcPTcxUuJdmv87znEr/x5jTn8n1Su9xccV/UX+DUGYgp2g244XLVl0iP5iM+crrss50vY/5
w3n+x5n104/CVhQzhbQGI5CEm8W6bYp4lKYxchPSVxKDbMDrKPynPu4vPRqTxZxJ92AsTtXwuUXR
3wR0sMzwZ0eAeiuCknjpuivRh52igHoQ3+PvfBtNF/tcICQz4Lw1BNZgXuILBHZUHhycU+gsdBWN
7kBrYJnkGPKuxsBhtvWlWeYAFECJxstf7IlwwthL1XWRun3brLBfWH7MXBDfqgtTXfl5n+zxMd0G
at5ZsTrZNZqnRCmcgaUztv3PpMptH9BqLGygZkwq68kXF0RiCpPOBt1K9vkE2syOXz11fwwZsTHa
iQ1aD3CDFNxwPyvY2SU7mwgJaI/s3xoFW1hMWh5mfuHvVHYReuNEL98da2+V0CDVcUpqYidDLog4
Z7Y3zt1OggMfZG66Z+Ee3UiqqYvZr2yhee40v7KTh85cbgsoY0MsndAGSk1WiIoCSn4wqWUKgHWb
tOo8WN1BhEmnS2AAMEkAvj5gcD+pJ4WepKAk9vrnJD8EiSh9eQtVGWbax9OKKELKFwnmDMLodMm+
ye1nFtD/zcOEJ+zguMvZfh3grP9BTW+jK9wAQknAKTP1UXF+SQhLNaZuWeOQrgWOxgebkLuvXTA4
11qBF2icaLVkSgXim12jlpRYQHCP0IwWjzJO23r7wPh012tbTf1Ikgqj6OLQIJW0JDWk0/i70nmk
6tefFsXdxznZtY1jxvunGa9kQSTJ5CRoUDxpXt6HCzNyF4pY7JiwivoA9LrZP1B9LJsOk84Q509Z
oLZwKSZiRcSLO/yxSiUh7iko116mEj525OAxZ+mA3BczsC20u0b60M/FTMyvKmP42SUdX1XmcTEi
D82GoUobT2b2OqXbQW9Qa8q2h0U0dSTOEQCtSO3gJaQYCCPcKs3Vqbs8KGZNYJEB2NcKCH+mw3K4
I0OG7i0YnDVSICK+OnyojD724yP98hj9eWoCWifb4YiUuZ3ry+Qv9xQAZqdadNRZKtn3faFsCVyY
4H66HvcBB9pGcncng+KPMKqvrYcWxbDR1jVaWXsQeIf84Pi9b4DyMSi6HNm5+uWmpDebvWvW8iLx
Hf2zEZQntczBzCOLhD351H6e9Uai8CVMlklaQmccwR7Pd6rn0dXLbe3JuHm/I3TUY4U8ls+hcFXo
AdYqNAYXIdy9W+VrtWRDpay3Wpx6E/m770SmimXJzJ/QcZg73U3FI+a1qzgP6fqhGtz2qfd2UU2I
bKW9C4ocOgr+GKK6KEB1FV3QmFkP5mL7KZNrpfZ9cgRaakRO0F6+3s+HNHL6H2ZeD/G+OmpVlAgu
Bl32u7bNFPSt8M+ut40vUa/o/ce1CIG4UzP7AmLQIgIl6TAPLuV0PUmWUgcusbnph8TV8ojF7jIW
vR3A89yBL8ONS50VWJuDIkKriVEiPgj6jqdpblImRMPF45Fl2YiurJuJwxJoqDpH7fYWRWp69t8k
lgj6CLXW5MnsjQ2PcviNNDyvCSHc6RzstCJxxIUd47nVnnU8DJVtDjuAD6N2VISNMYa7M3KDxq9a
DJ0INHjH7fmhK2I/WzTeZ6sJFj4Uftyawjij31/NgagAeJjsRCviNmw787ObSVmiS2DlE/8m6w/7
QyY8bP61vWbS44wFiBMaIxTIbsK+PrHWhC8fSDwp5+aCg1AypPnlhyzxaHugM65BPYa6uI9agNyD
NXV2mQcWWtO8+wJ417/XeWcgQO3jChdUx/opIB+TvxLio+DuG0wzlWR7G+MOKGTxnx7j7LbUHlXn
7Y15sOjayz4EYkoEQLPK8UNl6SL8ZGgU6nZXlpkQ/rMu4roU3A22cn7hplf8U3AVrjjTTOupmxkB
/1XBoveMJbl2Be/p0aIv/3787fA9Q/N6lN8UCqsOky9F9EaHfWIfVT/DWdD4Ak197VxrsXsyDMlC
h8Qll/oMmutXfTVCD1BKOXaqiscxXSw8hFIbDtUYfFWtjjtuoFxDDvzx3UP/I/s12ObfX7JcfGaq
yi29zhVGfAKcH5VKlTIctI5jGIOuCARuFN6UW67e64qpFlvwOHuvVsxg49tKMdIeUB1ljijt9aOX
N9wKEfZJ+MLNeKNlTMJgx5Q43IQSg3VSwRD883KVSpX7Ct5eH2NEB1hbp3OaI2oFzcDmeEqjHqSN
LEVsUyiQs1JIn8aN2MPIsNhmn5hvCD1nWlp0QEoEqe63tXQdF4j244rtF4HhH/DbPlmLOhrvIybo
zS5EU4w0yiUiC9Ft68I4WMIDU4aejcOxCcPse4c131GI1NX5cOFfuiu2+3GMCzB8qJ19Jf1rmV2j
Igjf/fbZ07cHTZFCH6gKXNW5sowkAOnN4gaV9KQr5kaS0Y0xrbnory4+zQpFRJEoqqAspn7IHu33
ncxCuy6NF51EKu+fLFwXIaZ7ytzUqzexREUuQIz4J/oEl0kZE6rpmAoPB06EUAMNGLZ+kmyxtB2X
vGSozNVmLMbPBB6jxxWboYefd9eBbcIsyKr/kACwMFqpbE0PrZ3w2UJT7kFhBCuz571dVz1hP8IM
VzWOfbgCfxD2PXhHdwcMxRL03s00HBeKCas0kVMmVFs8pC1I34yuu+2qzXYlnxLvSJyCiOVmgRnG
hSnTy0+ashpMTbJ9u520FXEw5xge3D1/T94REfRwxwzBN64VDjQ2dFuhxE5h1en/EqYYeCeZJd4r
ssany1UB0yV9Jr/Vpky67M7YX6mxED0tz19LQC3CioOTliBh+GB30SJslArozC0yPvZ8NhjGVj28
/TAObdThYarXiAFflyKYFlkNpxqcF7GRHBrduBj7QlzRPNLR2PLC7AAIqraryFq60jdQSuARhghP
K9nsPRIOQQhGKab7ZNPYLfNEk+OJh6LKprD2Erryz7zGVKqM6w+cwAj0QK46TiArNgj1ePWvV0Zd
TxLWmO5Z/GM6XkrOw8lC/syvk2HRCD1m08jmOrdJLWjIdthB6o1xtMOtjazLUtg7bvADr7OnO8ns
piezrWT8STawiIB+vavAzf7bwRn6NzlpeHc+JZhUoaC7Y49k/JoZCXcIglxBKWhePwwWC9LHZdtw
ELfcznPqNSa9guIHLD7YPcxTspyrQIZEUek4T5P/yidxDBcs836x96OFvkbFq9SXj5Croih7m9xU
3UxxST1/2Uzh7TqKd7H8mqM2wz7dTuYwApAjC/bU4hfuA+vQamWVooMc+TbIouHvWaqwvlzZ2FPv
vdICP6gRNhP1EtRdLm9Yy+TT4jWVJxLkwALj9BNC3SExBp+ZhLmfmDD1rpX4mmkpA4Ml34t8gi/2
wfZwdi6BwMu1DzdaLw816nLtMLv54KQxUFUFKdxn2/m5jDyjroRUimU4MkBFELl+VC4c2t9D0ccL
jN4jO42RC2lc0X4Tt8SlRF3dn0FNhNT/aeXj6e/rtjQWOO70tHrBG4tQ/8RLeJqdWtcKrgvlG4O9
RY7DLCQV3dgQsIP5qv9hbpFPw8sxPWukNXcvP6Jd9XH4/36vKV4l9Qo7J0bokMM4MOBUjgV03Rm6
hTlV++FsdvnpOa2HDJYYNqux+RzFJbwl11EBkMFq1oVH/lBg63xEpfG7sJ+V5nICVsFPIxN1bM2w
KRO//9WBgvISyrDeFXCzyN0PE9Ou5eqALTahePfNJjswIoYuvx9tMH0W6mFIU9c/0yBVoqBatMo8
k+Zdafq9Q7RyAKDLHgbqlV8ElyNwwLU47lCwYio2ZBUonJ67pRNCSYDYr2urj6AgVLseOrFy4L+p
H3yuVta/ujTpvr333EMrjDztAH/RlDcKEH6KCgTgV2VLHLbBMOmZK/yrEkY5WKe+TYHZtbhYAsyn
8or5ywoL7T1Toundeuc1Lb/XK9RtmLiFYsJySflLSrHqm3LulL1D4JSbfweG3YHS/bylx/RyYXNZ
MCBJO0WKJd4yUPXYWBT//g8XEDu+xrfiTJ7vyjut0XYEe4MXi1TRtacWYEpzR92S4HhKzcA5pNCN
g5xkLMT2oZMtFyuRTt3RiwgZXcnnhIO4a7F1qQf9YKpobYOD2HGFo883xQdD/SyZl7OGHSVkjXIa
N1aTXlQFGShbeGFo9EyJupsQD+35HxXGWyYX7rH2so2XJ5jrLONirWW5P4MuScPPzCjjAr71gH35
G50UozeDX07FlyanQ4Q+UScdLF/9wpCxq5S8cJInaGDGxXZSXrW+eLuQZNWhGh64TgLK9f2xwE2v
+W4zEQChfT3gngds+0h1vlITJKu85UsVS/z3E+z/1WmUXlWRBEjiHg/LYIwR7wfm1Dqh97mx4jMu
SxUw6K0rrRyZwsfuurkmo6/vsAnLEv9y/p4uYPtRjDMqqCuDXonabCsOafEzQprMNm/Ummwu8vUn
AhoEE08K8dq+nys1S6sAt1DZAerBhYLTPKSlc9X7P6xkXVZ6yy5GlKclO0eMa7ae3b13axZUJePi
uUiFB8A8WOp/EiNvK6U5BV+qi2UrIyI2bArf5RxOttO+1YMwZOYQDtAt1MKhkIw3JasRFIvcoTCw
l0VMYpQb/eOj8HYBI0dtxtF8msUkSZMz79PeoJW+ybGoLq4HoyFxuyOfnZ4l3+S0Rqc+qHVXWRCw
9EFKM1intn8u3IuKNwADSxQPW+y3iqYSFUymM6jxyrA8OExw6+7l/Mgkm4rmAHXheV2aVmQM6uuy
Y8ly+/DaxiWr80AZ0jxniPeRVDaYftL7ePGbHo7wQ+iGiCaopLgm/cpJxak+Fz5FqBSeh1i9pC3D
p4I956lm7qLB6glxGDeDDESb2sOfBsM8vLOU9kYNaViuWHbGZjrRL3RHjYtLKV3s3A1yDooATQD7
KdSt5TNHNSA45djFlELiyJGUXA6sVEeNaDv524TsoFKV81OUa8CEoCJqeHJS5jLX/kkOaQJcptDG
5rRfZnLkZK7G1dGDAdxofzkWgkYBL+hK4dWU9cz++ygX1z9JAGBIenMLGwDNlyZ6iOPJxYfUELu6
/7bGFy2nHv8ktfgAHsiuML1RQpGCbEH+ngiEG/k/OVLDDjHpH77nWSzD3s5p08IVpvS8xCKs/TWL
cuviUIqHgnMN+++I/XkWZDMBFeLtv4rr8Ho3PHoDGVHAjyMOhTgfvxMQZCI18MZQnR8ZCWhMk6Lf
SYd2FqHOgPGYc+J7jJ93mcj+95FEt6KmNLFnxHg7OUwE/SFDb2gkyJ9/u/7NVIG+oDYdG23lm2sH
DOlD3teSppIltIM/FDASxFrHXPO/f0ClRZZ6QvSlHU/iPcuUAys4pmZdbbJj4/4X16mNga6oVpdh
pe4MeAcGeIZJ83/Rkug8MbDfhoSCelvD15Lib2Itp2cckBmdhdTqzuwoB8AF0UHRN8SDoOV3Lp/5
OpQTLYo3dzFSMd+WbbfcLq8ueGD8tw2yhDxx6cm99wP5Mrqt5b5mNQAcicMMXZKw43WmCAYuy/TH
+QB83Z54h8bN5wXItrzF3JiDcM1dXaWmlnjz8GCf+ugkZRmHl+JpJ8U3St/URJNhn1AqFVNG6zQI
8gtJGgC1VvQ4c2qmhjGWycpbS9Qj+5ePQ+l7nJ/sYauy3NfwyUWSkbkbV05k2qOYRzSiH7Fhkbsg
S3gP+qg21TvKjDxTuQC+ZENrsw0RRgM020vVSkHMpOrbfEWnCUhPJh2BPhtLfJsnu9YBmGmR8dx4
21qeKLKWRRYknOvNK72O3dOsbOgRW/Xg7e9glxge7NIibriTfSodVI4b6ZmY/PiezgKv2s35rLEx
FI3sO1HLthPL/XKuRCRa1RefE0WP4PMV8g8eR5qDU0EGPsxTQKUAWZ/bgWQqMROZ9mGBIVHLzWAc
7c4M2AG1IHdGyT7wlo0/uPTxixMSdMI/DJnXW+sJnH2Z9dg1i94B16YP/ZCyt8fe0KykZLBvuI+k
s+tnaAEbC05fHog32NJwtyQmxBQcgm+kSP3p1iDVEcbeJoggbyyiKUfjK3qtpzFKotPZShBnAHLk
h7Whf8yd8A8V39SoZdK0A1A/TiWPZzFm+Cjc7vfZempDqVW4DbGp71azL87Kf5Ri47Gl7L3vwspW
45KuSFNkG3537EBBoWoxotqB5bDr7y3qx/lBdehgLuDRtQ9jJCK8se0OaUikMH4hMA5WbSMWxHfC
hRZFS5sO92JjvDcbuel+sGjaAbBR9JAF3kTsEews63VFMC1xmyyA8ziLKHIqUItClY6p0KlGQSVy
c6yLorZxYnkPYDEI7Y6ogve1PE18xfhJCWivD7pD29vS5YLGJX0vlDMUu0feNmvvZzj9ztKmbAkg
57bd68LpZzrjnmEy557NWPZonwScdxaG0T0p9ltxqv0aOPgiJWoOTLtGGMHstFX6EUgfUx4FWT9p
9vkc0jzLHYBX97aKV1Q5erRm11DzwCdKwYYGocGqcUufw+uJf5ye58IH30lXj75KVeFUH5UTm0sI
2/QAN5MHlbdMsbiPWapwRWXSLiI0PMjHoEYhV2UoCBeydZ0dAiv98XJuuZDCDszme1/wTImd58w8
Yss/d46BnwQphTk/coTefzDHmlxqJuZMKjJc8MREhk1Q0yIRoV2uaEKzgJxoTUQdlWx057cgK/hC
tVbQ/R7duWjyULuJHgMm94h4YH3NOSdsxhLM+o2f2UMBs0isqgNNFIjXk4L59F9O25a5Jbd06fBC
HIwHTMy2P05fzWkYyiix71mGONsb16w9OjOOOWsoo3oPW2v+YQ4GSLkvTke7CqYHgYg83XvORFCR
q1W4g8mPt6ysbUo9/X+lynLA8dGTw5A9Q41bhqWmfdk5JG1DABNv+Myc5SjKx0QoJqrHhLtmG1ff
KPftR1wCivNJTQDtwKR0tXF5pEYi/nSgW5vtj1pdFaXivENDQ66bpY61/7WkIjPQboyKAoxUiWcD
201eblAQI33Bd+S4rj5Tfri/2FratQE0zZTD0Q0h8sENi/CTDZGvNh3FkeCkbGbAyXUKNuq316K5
vccrOY/lHrBX+Ce5+I0jfRMRuslF9M8RfV8XxYI9OfTKNg7+HPiTVAIo3DAIhm9xl+L4YzP0RafS
WS6d/RQx5+nzExuDO6DMYcE0+RUCGqSMFnWjvvnrW3RY2iTGomEX0rFZx+O7iDTN08Hvou4nTcUo
8MnG/8f8mBb7FP9MxW5PgBpb8lvm3UZj8Zeg3Aow62gFmsuxbWESgh3XqHMrInEO7WsyHwu7G36H
Dflim4BQ/8qIOIDLZU8tTJ+MRUzpZTrbsYVrrBw6gVuQINOm7AyyOka+dggVIB4LLSH31GDgMzR4
aD+zfgxgvbN9s9Yjw+0Um9xbk2IVxt7XrrExJLlBYYAsiieGWAYUWU3lZ5j6wtSKhP0kMQ/IKCUh
8144ly3fw6EASv55a8h1WHEo6om0Buwl1lUkw0lOEuhuweMwaDpO7YNqVEfOKYaghI6qlLxB8S9n
/LUGaym4A7nDgIjZzNMqernDb9YdeRxuqNiYPUiRqoto5EM7y/DFtRTHxxm7bg3iyOBngM/gKB9t
2wHXd999NR5XT3yRRSgsiOKm8HJH+MwSO9vEpAOeRQ88Jwl3G37uxU/WL1EuFWnfipAXBBGZY0rS
Pn9IY7/AjsXnJ9XWXZhFaFrq+OWT7olV++ycm9tTCD0/ruhFay5HK2RmMhAoH6eND/jP1U+iTFPT
uBQ/mAAyLqa+NY5a5Jgr5sXYEbp8b8WwB32xumLfJn99qVXAgWxikKdRJIK3lCPUw2Vmzs+zDKnU
1WnmnKK4gtRAGzFn28ap1fw2NA93Yd/I6EFybtqbAaQY1WjDc9QFBA1w9D28ZxlpPLYD2Op7K8Se
zGCenf0gilwgGUBhMj/xY5r5iaYURbwP3J0DICXvFTfnVxlj5r8/l1oc9+C1G8anQkSWA0bjFa3z
s++p0nQpwHWWxpQtCQD0eW6AfK0SNALK5UPwTVQIXwEkiXcwScgFO6LBPcV2TyJCu5eqhC14pi+5
MmvsQOTJkhW77BTMPReppLz6PZZY56LF9KdDJq1yCf/Rw9dY/htZzG1//MJujDk3XTH/h/veEjSd
26GQHOncfPVAHjZyl48hVj9/+jhOSzF1UWCo9sohXQTWpxBnl4MdxLg8T8Z6UMSQveOUbkiv0WvE
NJt7Koj+qSuqYxTr47GT19Zwdw+yGyL7DYILZNV9SO1PawObBF8z5zPfutxxc0E3ZqxUp/nNpeFF
HhKiUnLhDCN8+t0mWTdrNO7/2QCDqWX2fYTv/O5Yw5uLlwDLKhDwsjekvkFnH7MDqHfgVQ996qqK
6siH85zaL0ILZbCWkUPJue8VeA4I/F+jFjW1hNSRfHziG4ZvrQdlGUbI6NJTSHGH6+RSE7D9eJFz
pMBO50bG9JK5R7U95JEeyyW5DUu4cDxLZ0cLzi4ygLobqzsOoA+Bs77Itv/c23qoHrXzWo0Yt7xU
BdmBKvAkpmBLSefKLDaC0Aiat4yNMIC+jr6to7h+uWHiPYo3seZwe+6LnxiDhLOvaF9dJF8zJLki
tTVQkjEUdPqJz9QhOqMo6zn8kf8rq540PYF2sK/6rKexj2A2cfIF5D2fadSbYZrnqOXWiAumBc3B
n2aLUtu/kSl3uyF8wh37I17pcBjV7qQGUjSLaThoGSiZ+gkUtXSuBlK/8m6JUaB/P7DUz8gGlQZX
Lt6SoA3lI3o96FWIid+Aq8cosvLDV6cOEZEHVRHwHxYOugx4J8DXDm5TEl4vm+UMjSJcmmC2ealq
xImKyO5uZqIOBSgtOmVxhpCRD+Q9PkDZtY3xakXxBN+BrpTA3jQKfXH8FNM9NQP2HJJTKOi6OjAy
ttHKlFm9CTXoBjHB+/M8fg70AJNzaR8puc6kyrebzx/fgWAAKTFpO85/6FnTcEy7Bh+b22tHTMy3
5JltOQmZoJM5KS9Vq1g3FCJPQWwC3jb6dyyyFHlft5yrXFardnxjzjIVNiLZEfBSh/OnnA+vHlXg
yIsPpsfSVqgV7lqukCzE7gK4YnjjmOZfYTxJtpYjFgWq5CbSf6oox7ldf8B8QHbOrGNVUzJC3lhj
jeewoH95Zm8U+OpuMAC/s5+RF8zN51KggXMO0FhGVk/cqKlevvWQbsS0p9Ey5TFPNhsQJmqdbUBu
iY9z2bUfzTsNQnW/haNZB1Ixh6qT+JANsUgEK6kdVhm/6QMLLfPILTq4WDIo3BA8u+c+KprQemer
4D0kZjcp4jGI/Fa7vqGM+dNCIJDEkS0cx0POpBmZjkn5LAoZ/BHel1l2SvVuwSKHJgmTwlM0TOaE
JhqiGnvqZxAhBecnbbNGcquB1KqPmjsqifva0ZDGmhUkoW16mxwwwOqalPXHjT4A+tf84EceU2Y2
A2SME93gkSXspu+eiPqPxqBu2AJx6mcUA07wFkwNjP4rKDENg87F+jcQNdMICkQ+OHWN64Z3BL9C
uYZsN7XLf77G+R+pjZ5lK3ABLsX0cN/ifuR+da8Zi35IMvHleBlc10dRPYjQgxFxulcbMushcTcN
y/BeyeRI15Vp7OL9/ZUIgd/f0DRL3qt3+JY3BlIVLyzQ1Ltf4QbQ/a5NG4MSkhZHbaaiTQ0KNrMf
f+txs0sm+4yuuS7NH1eTsIRD6iIGTfSRhLxz3owY2LKdNvWhb0g5JCFZMxJF/qXe6N5jalYcJjbu
eOJU2YcNqpbcb8MyxjWFS8bMiG8T6U/qtxGJUODJZwJHtOKZhGhyrfjS0Ef1CJFkulCD0x4GsvJD
BgL/nKQW+3lxdtxswsU/3/i/8nQMrXmfu/Y4V0VWrXaTnxo6Y43MDMcLicmcCnkFSKIr+pNEm8yt
MXUg/6BFiYg7R7fm1w+AJnrdYRZDk2DtxU+Aj/Nu+ZCGwhNIMg7CEAggL85ILRHuzkWp2UIY8PzT
okAQT9YJvn4OuKeDziAGcLo1cpEzF6lnyhlK+wz1cwvDE3ewYvQpjEo4KA4vlUjIXhCH24GBm9+O
SaORUsqNcw17TovKmP+VH/u3mrzpSgrY5aCgz5tPFg015T1U+I2vecPcgN351u8jErsAshbKINR9
fVQQZosDl/+vp60gJpJMCujtxDO7/tZM/rNiBDAJT10FSc9XBPwx+TMLc1SRBgMYlxWJB2t+sY1E
MPlBckVkSgm6AclK4MCZkQhhUbi0rqTPXeJwFdQV2rh701PIS1Cu34Wagl/ZHAGbgYxxFd988kox
ydK1PtFbqZJqRx+LG6hJSYnqxp62WLvMugBtSarixTptPThHOdiGH7PguKWgCivEX0bYtc+QYxZR
lyCQb9jhCXr7XPE942S1E9tspIjKnnkkwVWFArrHKsIENxBlVT3f26B7ldTya8Di4ZhpMaDPhM0F
BlSLu/3idRY5BHW3JxGVa6+2f+vERwWs5j4M5xDhRLn/FvCMg2rpwQXNf8BsuE3WHtH9kX9/i4jI
gAiCAR5pxTAyx/gTL4nqLXVFqzmzeQXnztPtboEW2OsqVbRwnh/iYRxO3hCrH822Up2ewg9pW6P6
GEhWlhbpQ+YSholqBjRgsXCXNyKq2bcHwanBFLZOzLuqOo01W1Zn54hT2KlrdzfxNYGY09YxomOl
fI4LXqmUaW9YeiVig3wphYiJjGnEpKQvaj8FsrBDqW4eXG5g+Qf+NFXRwdAtpnOXy/TUuW8K5Qeh
YLehHVhZdsMMTyAJO0aUNoo31rkAWD9loOgVsttCtEvrSTNvuLPQjIN4cumo1tYsQkpaDg4VNEEj
rjAI/VaVdrMfnGsMX0U9k+na6T6KwY7MyE5sAFFv+iHzHTIvwozer/itd98z4ePA3CCMCT8bFmaV
VuSkuqKJsmBO0dcoOgLaa/WPL4UsS492qwmkX0uaUYSlQijDc9pbh22LInKZ2QaeOUleR6qm3Bli
m5Kx2Z5LiC5m3W4pGzJXE9RR/g4wwmMRRpsGheUDVwbfpDBjWUEwYxj0ymsd/oi+LRZvwQlwUcL0
ePR94Kw8anHihmdoWD/oesYu/Fh57VHf3Gp/QW0b5w9uaeWZKjmrFVIWfKEtXLtnFtE3IyYFwoOZ
KKj/b4QlNrJPvcHIUF+EFCxkkAsX1o+/LaPsNegHULtfYItQ84bFz/u0P3zvlQ6PPoXk104zCbja
oYvT7EajEcgHuIkCmIg9A8sZKDHmCaYrcYqCqofJl8o/GEXolPMy6jSoXOJWEP9b2oxYCyKChzYV
3Zl+rFFJNl15exObQZeYLMqGL4c1rwjI1BfIVdNwI9U+VHWjb1cGbcQD7hAZKeGvITCu22UMPgYr
za7i874nkgJfNIsfKy89tY9vo/60AXFsl4r1J3DOLjKwesdVa+r8I+kYb2xGAUIx0HbbDKFonImv
vuLjog2oz2kNjBlxrqHt//4+yG4MQYvdgroraD6Y0ok4XqikaNNbOEzzQkVsg2zheDH+t53Mw132
ACmXuXvCRyLHNV1X/ih9ybAdZ0uWsRKL+UNvPNfy0qZuF6Fy+tjOuQKhhhA7hjggEYEkJU1yLm2o
UfbrvstYmReamjei/8hyorWrUXlrY7GkaZCp/HpjO1GGZge598tDioHQqIb4XFYETSyYVwx6AuZU
UY8x0hmjNh8WOx9S5gERdxGTmQGL5kLLnAn0dMhpXTb3zHHm6bukdiUHtDAe8m3Aw8yXrkX/Tjiu
GMGIxx7pQHi1+HTe9gbJS+s4OvBNszbfqT+b/Z8iNWPnVXDpfL6N3CWZLLzT9dp4OPlly95mOlcA
VUd/hF4+fjNSdHORHoK6w8QrUnBc0IGMdw5ufI9C0Nw3JN0D2Fk5zCX2AlQRAMQNew6nI36qz9wX
toc2pEQs6p+V9s4v4Bf7hwFKgjD/Aj+NT5vdCb2pNVAG5+anfTx1Vkb14rP8VaVP/8rDwZSLGxrF
9uFvmU7bZUvl53XCLPmnrVvHiQBaWW6FPKdR7IL4XP/FX5ltA4BgYaJWTspQcDRSl+/ZxKa9SacY
nPPPXCU+6OkQQR+GOGtsHJFVdyl837CKOJ+WpqQqnvgIeohr9a7urtUuEKc7po1SiBAEmnBtV3b6
JKWyfPPjvqNMyTb8fX6H9elfm2xKwsp48dfd65GUFy6Kg2dAeGcCI0eYnz+fc21bqbnFpxFjikJU
g42/WhlveRJfF8XTg0W6nCqf2eS+zXalL5J75pbS+EQnVZ6B5/agrRlP2nYdqy382kR8I4+xBliY
cYAhkGb1FGj48hCqX8A25tubjECcm/gcqVvucU3zhuzW5clomEFxBnkw/0XECGw3435QEJ/0GXf6
RVqaEhy5UwQ+ys6WESCOaso0VTJB42KOxwDx5ryMQcIxuZlFT3O4qb2VeZ2l05jqxP4L2TKCSb5/
1QznuBUEOO9Ywb8Xo+0phPVFDhhQWFGBeRe8tg07sUmKz+TH7kHPRHdb1RlNM3U8ThqQH5q+1KAR
DvPZo9zrQTagkBnz4uOI/XIF0k8msSTzCXvz/LovXLPMqvChihtWQIntUOoLZOCi4B87n1z3OdBO
53WSYPnkpWb/pHH2bSohWfJuxHCdJdAM7FmeaN40KPala106GH6BrhBo4lUr68MeMQPQL+AtVrwL
h7jyPvQd3rg0NXgKXGHBv0tCTEwWcZoqgrgW00xoZSnuuiY+H2en7UWFPsTGuuVXu0KN7C7l8e4l
QrFXh4nsb603+te9umkGGT7jp2HHU88PCbvnbSsz23MLMlmXx0senFwcl8qYhvl1n+WgJIqzvF8I
LhwHmsEaAgC6c9mGrDn0mj5v1MPXwi8Ul2L7n+q3bO0H/auFelnMCJfMfQzbAUVuRLquAs/GQFnW
jzGEN8VqFe7mKm4ndzh+q8Rel1Lgg4lO9/1/gUubkiUCOmcPmQ50tBKt6RgK9j1Q7uniwFUaVaDt
OV7nGqDGeDYX/5Hoyh//eSg4mcxxBmlzjqbLe6NlpLY4guz3/W1AIqJP+AGBTejxqJo6TFj3Wxa5
eIBi584yIzTSAp1uSHT6fPWdzTxGaWf3OWdLisWl8CneyvnTOCqRGsQrNr8WR+YSC+GFR7kwKGAL
FmtH32g3vGKqN2N69kInNCds8gegkGxmmu+/Cv0Qf7HHbdO142CscoyeVjOx5m2KacO3lnHij9Rs
96UYA8oilMd7MFQSKryl1UFYWx758AfKcKzIq/wpuMNxE4jaJWSolDa6q6oNY2igj/9BEAZmd0mm
WsMzsKdSte8aN9TtHeLsE2Ux17JOIVLsSjjks9CNHcEJYwrpKU+S0aA2fyRG2R9lCLL9uo1c9fiE
JzfRDgbvOM42x0Vk+AihHlZFZXfc3sgafhraW2uLOBjSyTDyQqLmvd6x2D0NISCb43CBaX3CNGDI
ULuTZqII3+26cefrPMhmur56DY4+Dub2/1gK+vHThpGGfgk6qYgVucja5Xa/ytHq0Rv05CMoDRvB
8gRZ1xVIKttgOihvKcUrpMMSAlK5lmwR0ULrS5zA7oPTRdUiqDOjGa+4Jyn4Bbv5Nh8jJ8e1y6Md
P3TY1S5QHgvUPxzBVJjpvPaX1Ti++/g6vgvMM9Mtt0vNCfCN1soXCJGHWgxlKj2J7rudZz0JkIFH
polD1U/dVIVubccABYjvlU6gFD7LzbjPwtfVmH8BpP26hz9PiNdrJ5bEa4IOL0g1P1UST+933YI/
rhZCC+CZZMi8TX/KIqdXdFJPNzWXgHc8erRfVmqCD2rZxfwbDfOPBSN2BN7S3YkP0WMNiV1VjZN/
Rd+OAS0TN1rtpvFV70176lVemilgYeJIpwaaseHllN1CQA1/MLoV1RrHrzOIR3TpmGs9qVNnGccC
s/ynNF3YfISHpmnhYCtMEQB0b3K9t/P8xX2ZLMgMAMYPNInL9JatcoM026y70Svz/zbXg0cXgrq4
zzejeIU3VNhrEEVBDzidhJY6rey9Fdm5xoLsWFFKF8wQ1NDvk+LKisROCUqSreh6ST8gsepo8Spi
uQWthm5nlo/9n+iMPShCSDCLzEEreThhiFUh6+8k1elyxzrQDgete59xD94zrD6uLnsp0CVCYdfc
Lr3i+NZwrFCK8N+PkCCAZMu7PieNoI5InBvrBJsC0y2xXJen8GIV64x1zdRgPhAuCXYO3v0HTxhl
GNY7u4CAT95JNDk4Up3IeePeRw06Ghf4hem3y6A7C7U8flSIL2SGSFPf7rhAbXBKIKB3a5LCU2e+
lRPCbi3jjA7TKBP22Hy0rENnp3j8Azx3mEey/Z3FpD6DKTIFGewTics2NyK3nJU9JJpt6jndyQoh
HPepPq3UURfSaQUqBpiM9ZHH/zOgn04zH3MqIeRoukF8VQ5X/dPFLRBt2Jo4Bj9p05sJ/E6lBnPj
KLMsq0UGxbuaouWUDhGRrzUB4WF6dakkfgmcvz+GdZtAGywKS2AjGPPX59PyN4u59ysLbBKjgyGY
nXeqorUwt6hdsFn9io6aOpsB+eV8cE/hu5Ftvk18vFwvYI+OrkwxXlB4kMwPLbXJ9niMuD34A/Tp
p8NvMnXjjocHE73cZ00AJbyGTgguDQthx14QbGb+YpxyA8ba4wgVrFJbhbFVVZibQMrPlTWKWkCk
18LQVEz+iR4qkOCHfKswScZQNovLZmtViFeKqYkzb28zfAx+B/ARmMQKa/wr1PJGHOQ85yseyY2Q
1ercXKQwcch5pqE20NfIA2tvSSE/gI5f/nDBqxtthGElI0T9gIuE1Pw7tqpFH3Uv9U0ggJ0KC8Nz
hOVh45kocJxgsKCnw/qvxpq6VpmbOUaUfpIjcf0RjaQfxWY3WeYmq5khkg7qJkUOMzhumugem9Mi
GOJJL5PJOmRov/BeoyK5BJtlk0gpdQLXI2cyLq0/yolz3cKgvPGyEjvuFwlvlprpGUVmunMQeVI7
7J6Lk57MHjLPLHkXi9WI/wTsVmS/4X5N3V2ldFDDTkg4YUg4zYMEj7Hrgw0Ut22V5oUake5ahEqE
FMRl0gYsy+BWGl8KZsJpG9Ix72P0pvdqex/99EYcMnLW3x5UqTQnTNd5kCP/e5vM2J8LnLjENM90
8dbqlUzWK18tfkDpaQ38tLaRXfDxwU6JlC9qfxo88Zjmu9+uFwYxsHHCFQs1eU4w+SM2PxFhiewk
RCPfDhP8EzN5OY0uSCKkjTRVkhvTBuxCepItiW7rRgOfChtJiJgTuP8NUxydU4cA61IihmBG9sJJ
0wQNlP6M56WH05+KQ4bGoD9MsvZ4yTJHXnV0M0CHddDlHGsnW/GdLR5rvDEzO7RJKVJ/btSmcTQS
51R3pjHc09u40RFzfwRfqCEhFONYuuSmhl8qkULaPfqYQjRCI+3zaiftB/u2075TIsbny3uS6oeD
eSiGxveVsD5/0qbggvBvbNujTXdKo6atelBoS+GCE4I/S5Qge21k87WgbW3YXyD+N5UoE+NvvWfL
wTaayl47CA2r9H9JeF45el9LyNsYQKQEfQEg/Wxhr129EKazgCUmjQdcxX5TsxYYU1kgLuje+LcZ
Xa3WITZZ+9y/YhkZn0qULIOV7vy8pL23Vo2vKcKgoSCd8duwEKkxY02CvSknuQbL6RuIhPm/Myuo
hLJdr1LtHSRWrEHeYULNN5jm9uUsgmByGjRVKV1ckeXfG+ix+as09GB7cfI8qXPz31C8SQiiLCyZ
9LcORA56y2Ux3uXznFcCxZfbW4uLZVOw+CDgHDRNLKEJzo33nb+QaWgMjIJg4m4gKNXx4eYyQHT2
DF8MgyFNDXPKxarAaUBNAURSJVNUMTfsiBsQf45y+xVSErS72VIEpiW5VqmswuhNVvXMfutBdZB9
/4UJIHIUI6JUWyeLHwRSeeaNeHwUU0QA9o7TRNjgYSisV21FzCZo8D0NWotpfPEDS2lrrBpEZOrt
45qafPIBEVNEuwY32/HlJeKqhOYTOmNgU9cdYsKUWk0pdswa6fEtBOsTYHXmJ5To+bYqrYRDKquc
tKcePsBp/x8TcoZ+jogUM0AcwWJKXTu+OF8n2qM+iK/UrojImLahOWcJcotrHyrVJLh0II+8+Hcw
PwzZbEMyA+FWy5/NtD/lgfLVVo0D9xn3KovnAZj45dxdmtWUGdC9/UbXqE39VZsmmM9UdHaBwViX
oNOdLeN+fiW51ZEmzAHDPBOklVmPmdPXg43iN/XwfabeuQSQ2yA7RV80+w97ZLx7Z3cYh4d0rmHl
SYp1YOkBCoothaFZhripiTTjURPQDohAPGCcY8Fdq/yhcMTmEbYGrWDmKwrEvfDykUccR8zNZyGR
f0tQFe+pxkbe0KvTuntP5hBrg3UKju6RWJAvL3DNlD8lO7jrPl1sQ1Eh2Sh4rGsrBIMAXx5fg9ju
JjMHwTK4z+jVwK1CfvaR12q322gBVqMJ0OcTW0OH32kxPfwyaq6qA/OXpEXukmBTiLPiJcZ4A71K
2k8UiDps8bOo8FceZWWT3KZ0UXlBzaUoLOfp2i7SQNRK9Tr5HXrBJa2AHuJgRlQnONBNf6Yguffn
eSl+Asa5wW1BN6Xpu9+/4CLdcpyt7EP8e8cqddYCkYg5eqBPR2fQeqmSoLpfhVTDw+uSLPRZQHTQ
gPkYwFlNuNYEHwR5j2ko2yR/Y1cxV7a0euxzdk9RVzuDSq5xI4F5HVCSyuiKydxm4BhxaItsRNIt
bKIlKIJFzWxa/gC+wjG+MtRmN+AZAvTbWb3eSYZvpOui8KNpwXISPxXuNvRrtkYT5SrXCEURlCW3
uHC/3MJkcGbQNy/BItzJ93c4Xv/6rZmrpUmpeVNbP6yKae98s9we9Qk0E3Ku+bIWSSEW4JFPf81D
tDBF7Pe3U2W4SKjUgIRepfrEkmI5itL0DfkZ11fTCvHO7o/rD7uu5MZWp2nSRjfi/H5vhuG3GbfT
igPv/odos8xKuf8UB8Hf4u8p9pk+r63x0AS904j0ck85oiCeLiC2KguxTGSnCVNmYf5W0/3aArPv
QKGS0zz41pNja/yDC2DFAP/3c4diVuxDOU/Evc0TYBIDlp+3Me1JuBkKZy5jD10q84HJ2HW7Wrqe
7xjLs04ndhLOTywCalGJa9144jOmNBGbePCrrgX/Jw/OpLzgtVxPgFMZu3HsuONhNBw4pXGimCfO
C8ZQkhVH8wzFhoSf25YKr1JvmKmjRUnWfIQOEKfwetyv5tSC23nKcPjMRQyHEStPSo/VVb5O1hVN
WHkuZSmjntb9GKoEV8OtCQ11iHgNdE2Y3ScVI2I3O+YBpNvFC8UnGB3YaNNyj9rFOtxkt7eCo4Fr
JwOUh7DGc9SGcPTQJGcbZEx/cLDmItTzzocgljrwOjt7E5xbvPexGyMu4+GvJECb6iiBg8VPKpXg
ZDHcydMr3Ly7dhSsIh0dmbD780Blfh97np/4yNnX1pGIRDj6aX6RmbQM4A9JltuhioBzJDLMyOoZ
3MLNNnfFZ0/CnteYa7BQJo6iiegobHzP6oRVuaAVWkzlveav2Yaxk4OiRg26aYbjzUnEDVvbXyDE
mdA12dmEemz9ukSNoL/0YDVQ7YV+HtjnbSWtrCqriBLUmDO+LnaABdvC8JQ/t3GPfd8AQ95kqT5y
0cVcmhXE3mJU+PyhaCgnOdDfH4XhZVFta4icV086+35vzxUpLqVvIMi1OpjPgE2rtOmc72iw7o69
oWgQyvgejezO2P156nomgpQgHdb1zhm5IHEI0IdVqcOt9Qpyq3Et8V3FKi2epNSbCwygHsY/zpwG
dH0+sKWm8lP/r97ccJVHFZ4z8NbRIQCQyv6f48D3/gBy3omd3Kxv8nvTy69H6Z9uejjRvvtr50ic
OgYYtP3y/xwlcoKldp8tbVFB1+vSJgbjkmSiY6MYCMfeH0u7Obotzj2oFo6UJtCdYOsJHD3mocvY
MVtks9oC+/7b5umA3QdoxYUsSOxjJIzm/Zd4por/Qb54MIyVKUWFCKJAmqCK3XfFsk2ofxkZekKr
Pb6HGfNG/7SrOJD5NSkfzKRhbDVVeOU6RX4cGwcOpfeDgIVpjkA6a64K46maO0YGzQAO+EWLOOKL
Dg0tR/7mmFFInS3ziqE7o79YKbjkPSkLj/irU8QR4c85Te6ra+jHRW2uAAeYD9tm5apoMuMoLyWg
9zI4pB1pLztKNqnHSsR/5a7aVtfeNCliK+erCTEezGJTOnPjXfQLNfyCl146Ey+JKaqEzX2SABn4
HMFmt4v5cF6isfh+XjbsOGQjHl4II3qiHTT+ffqKBQMYaPjNvoSsOgYsauCg1Cv6YUmnt2i+ccA9
JyvcOpy+YACGCkgU8d2v5oL5zUkEAygd9HVkPxBxrSiGo5W4uYzFX+EIE3S6/Qvr79W6B449IfUM
KxwOnxXuSMAsezdOdXstsvtsgaqAC8CY9ApBNOJtTciKTmStkz8ZYyg4RV0FrcWN+xYSpNQZnOPR
EvNHl5EVvMFYbZe24J/97llViQHyvtzySBnaUNH/7uzCUEDS4tiDSM7CmZkjkF+2HjoX/2LLevYT
YKTGShHSSe87kqhLlBqvoo0g9FmSDP1AXMKwj4OvVPjUtuvbUJDgsj9JPGvLCoWKTp9+v5eOK4ax
c5XRVchLXTemiLj/RHoNbdRPZAI0oUYHeHD2VRYoPw2vF4/UmgHmhLp6C5EiTYZZgwENd4Ask2pQ
2ywQulSRDgeak/VkiaGNYpSKbGleSuUCCetMMrTTFKheDugKSCs3dmGJhdThHoEzOOk89jlYTcVW
wi5fuRczJ0rQSJ+QTH7AkMaC9pw91z0PLrQu4xUq/cbx6SOQCGGdoTu9dI2Agy3XoIkI8JsmlfQ/
Zjd2x/LU3w2K0aRlhaGk9C3mhP3rf+cWeUPnAh7U3LhlAe/Cgvcf0J8XuQJBrryfFfJRqDKETos0
mTFYtOXWeOTdElxbrkFA/7y8GAIoFY7/hhSAi5fyoqFetnjPoMSIiOr/07GbN/+ESaixwdlzmVpn
/8BqMArwuSFYaUFBeRX9iXQpweZtOVDgmZfVsYaSswCmG0DXc1yyi4JCYp5rlrQEPGJC3Mi8A6JL
qf3RQdAVwsK5fJHux/2ZWLs7JvIpseR/qTe+ZQDc76TJMg0qAu/omCtx9fyaZRsn2L0LKVhNq7/3
MrxepoErA5dsk7PLHDCvRBCZrSMCbDPV5IjBxge4hnXq2sVkt122J8MmNKdx3AatCR+VBfH1JJES
+Zu+IIY/hs1u+JYSwlUnhdrskbQt3JutzGIewkQ8zpVO/jhEu2H9qfXpoT90gVj977qASNwvK/W+
H4q4tV4TSoLbAz5clo79M9602vjIa3oTlSrNzBuvy0NMb4VvGlMqIozRcUGHZBXB9XtVEhTobSiy
iOkZbEKGl1TTfw9dmAHvDf+/RjyXOUeNbqUnf25BQ0xnYe+/yVJqUGZN13aR6Dryhu5MOC1C92Kr
2vN9Ban3YHBpzA9jeTb9ZXshHVr2KhLY9jbb0d8QdX/h0I8CDFcJEzo7PsX3sMGtA29rFpwevn5/
ptQZa704s67qPBoSx07wuRopNyuE/2/XVBRi8QZycRi0I7crLmA4BoOjJUI2VEJTTwCNsY+Zi3b0
yLfY3J2rY4sWx7UFaDnQbKbmCypsCvOewbrGL7ShLC43v3ivB1m/Cqjd9xCZyC65BEHMnG1632NH
IelhRpeByXpu253egI3Lwibudk/G44nddI7Ux40JwkclYxTkLzfHZs5rVYdQgJbkpkpLg2QVWYDe
2AZW1idyjgBJ91bD88XQguhKsR8ywnoi+B5I+wAzbgvzTL35qVBWyglbK+szIco5qkouMD5eZXMI
q2fdwg19xY8/MNj0Xlo8zSQkYQUQpfE0u7Vm/PVtdwI4lmL7+O6lrcIdQJ6zzbf9U0kFGl+66MQd
iDcwHWSLarjoBYA5yS07NBUObc7PIoCa+V87v5kXnGXv0qXXuBpZ2bb1mcb//gd3kzXUELChLDej
gndiKtxlmjvB9WCiGPG98lmfhr+UYf9XTwtcqgHQ56mDyeBlc/+nEfJzJ/Uu/z1vxusACVi4zAKz
HOupboLltBHPK/RBK3W8nwUClK1dhAU9rIj5vVNbohQIk/dxLZClOFft/FMKp9ZvHldhOEYJWjyZ
SLXn4nRS0sFYir6vGJazszBWl+jPtvQ9+iwkK38jX8jXU5oi2Yxla+b0IhzQcFWsFS2iUuFoQXdx
j5dcrRS0a95OHaUgP99ezKqP7OZsT0PZk8vyMWTTx+2akeQZODpHoIpHV8F50bVuSxd1k2yQTkak
k7TT0hfMGKcKnYBCPUue7v93eAhfOLPHFcchQqLOfE4jEgG1160ZwLdrNm3hKaUesT2e5u/ItApD
YwuQCkoelKTfRI/nAVH+Et/T5DuB3jI232eGjEkBlB3HdezX2ZHc9KnmM/RZD0Ns5k5S5BJ4ZmJV
KIE3zYU+WGOO4ALtRItErOBYUezmke02iso3FXnDURQgMLUr5o7cov/fZMBPIZOF+Las44NsGKqy
OYDHf0EA9RYQkb8/KlIR9ItHiPlKHiE/pfewbRFnsrDvD7UJzhiIKT3Wha3G9eIi4ab1mLlDyhWz
KbWVW5So94yACfiP7LtntCEgPiL1lVoeGyZHFYTifTsKQjCVa5Q6KgOzYaHmHED5nCwuzb0HEYKB
+3Fd/06qJIsbYCrga3A/I1BNhDHxknS8mmLONPRCxxJj9FuyFzmhS04tr7QVHxGlHBcNOSH7kVS0
lgK4biM6qXvgRK3m/MxQunrTzEjx1MhzJy6pHt6x60kh3aCM8VwTxvrZFXJZxcno/gFQtQ97u3/Y
mcWJUTeYzr6q7xBRuE1KEN+Fq72cn+qru7iU9g2pmMfBYygyYh+Gbe782gLtXSF5EcgYNyR6oMMe
8D7NKo8D3f/DIFYI3REooiiIdr3pcGYrTdtJV4K4fOkxHACL/I1PR9dXfsYrIWSu3GREvd5wbMJB
vv8k7yWMxVYkrgS5jE5aVALQYR9C8PcldDXeplxWB4sVUEawYv8o2oQLrIWUuzKPMmhvBCznghmj
rXbWqQtNiJEdMHwZ9Rw4ekybEXoEYssmKaM8upK6+Pr8Flr0T4DOlioJmdEHuPbQuF4FZNsEYOvA
o5Y6DkS3xBj7qRDcxgcFpeS7LyqmVF5S/HcbW13Rde/7N1z+EyLMRaHRYJ0yuw9OPc/TdDIb28DR
I1WVzU9GHKKGJv8QsHgwuAY7HePo9feZtWflj6CUmgMIC4DtdLFsGrrkV3E/JZj+batKvEJhUllV
x4dzPt01e+yzCM7HJh7Uqi8GQJZaZVaY4GXNlTgvTvLB9uwB8tNF6B7nK9HFn6bOqG1XuKDiTKg+
EZcUOCJsss8hqQfVv5OHGl5J9XCPJChAxRVm9O/SMcV658RVS7NgEslcduhT0Wl6KFWWq8F9h6Fz
782yJheUdP3N0G43k0CoV+Uj+U+DIgWm0ItR6s/H/PquOm7kBGZ4tpbiX5SAUgd7ksvBpamuR5Nw
4X2rK7L+Ojg5NPs2wHX1y5NmFnOp5xKX27dekChI2jDiJ49Z7cIR3lRf2IXlTrqYw8SRQqYrZlW7
XWevOVwJ65B6hGHfM9b373OnU/4rAGH5H1RIskS1We9vSmPii34ePPuJXl3Vb2j0ITnHuhECJbvL
tgRaORHYlkak5RChgoKuaDCa6P+57DN5bBThNdTYvpdUoTJ5Yy+CsNypqqYHls9UtYLgU6QQCJlh
yl11ySoPzpzDsRXA0MGaYOZ50CTYqM3kuldPmwXGTtlJl9/yx4eW4Q821oz8SXd/xyjJSnlTz0Pg
ymqsW5bFP7DpxL3DWP43tU6BEG6GTHuFteebltkK2Kqn58/UHFbW0vQUspzjXWubJ7EBoxMI27Iu
IS5uFCWkWbECnrsvLTTFRgg/SHN43jLNd5UrAsEYezT1bwIrkHZRh7TgsarxIFrCOm4UlJEsTmyQ
YIZh7V1i8dL5d6xbsesYDUT4BosqbvuVCXq9EvBj8+QNRyOaiSzRQNm/uuY1dgONipgLxoMoXR6G
pSyfTB3OhOE5X6PCDrra3XocdY1VqQWttIsJcyknkFt1qvF4FmI+qOLDbDXl+8VF5Co81MUbz/V/
hXnHUtPhhszcv4ippHdoZmjqsIzihq8slBkIiThonhw/jhd3h46D3D2KzEsUokjK8FukRSPbPd4q
D1zc7cuQLZU24pL48h0Wxl545xOjllu5IXHllI1oWibrnK2cKjmRNsuu94jR3oUQiRYjbdd12Eus
tpBmPGrqP+CV6SZ2J4n/6Bu+XtKpLoJaxFrrH8FtK1mxN9FbwVTk4a0Dhsnaxi7fq3t/dKN/Lyhx
VUByf9iIAzig3bdUAa5DueX6GM/FFV6Z4qftYwOHWDzvNOXAQXol9S1Cn5Brrk75Dmel7HAwVovM
QroCcHjA+YAJZv5Va8H2kJlIv+3pwd1xndSmgCEE/DlztsMy7jHRwcLORVvw28puiiBqCm8+hqyh
+Ta11m88OkEIjwAjRlIwts3QTRKaKaTTCe1H4W/pWPLiQRenIgkU0qaCnW/IstgReG0t/oZgXLjh
bksFzl2Lgn8uxhKLic2wEg2/GkRvCeTnUZNluA2vJMcmoISEAi9iXU8PrU4/VZMhQHBd3ffCpD+I
UXtePlqDfkoslssuWIq846cbZs8vALY4HBgZS5WzP/8unY6o5o8wGQdJ8AebwGapHKwZVhDOk8Zl
KkbU5UPbna8vAaOe7GDy8RRi7xpQ80fesNCLVwfpk5NZ531/sCQL4r4WLis2OwWR1vTJ/Y+TUhUc
vJrCqMzxj5Jdzva5B/TMFmA7wR6pgML4PL4+cIQAV43JsEqvbiwc7PNxPGw6UfnPrmdQiXwuiJj+
IaKB4SLURMijvRHWnXUZyreGu4bN+9Se8K0b4+4v776qPzXsgG9bnQfWC6uSrat14PH9u0AKBVR5
KdO9noU9+r7tB/0KI9OdIXApQMN/YvG0ZIxzflvIyD7igJKk26H7uGBcEWp6fLPBDhuaWDwCTru7
fT+0s2gK+3I7XTSezBLynGrL/OffvYzDwXtwJY/K7eCA4gk3SrF1SmRJ6tHlqE0+0JIJU6jcEHXm
wO2aCdfu+PzhoOk8Yi710AcKLmNNMTzVm2/sY0ffzWFBmrP8hue57KZPfYIlp+MDs078mC+VlFlQ
MXV3Cd4u4qWPXXN3fXZqfjcrNx95VKhTwu/GnZ7GsCwh73ko4LEgbnakoCOae4ne8b3GFY2Xkwrq
P+5Bct01n6srZgnFx2AlsQHCBRC+BrF33o2+5me73e8Jze5TUhabwosc1YIG9aiycMK8hBFFXibE
/kNA++QMg1bS3RSxEE+4NfW4Jpil2KqzCJRR+1Ft6aESP8uT1g+gmEodqb2e+JJgJM7xzpMTuiau
qqthIy7WfFFKRSWwMylXAc0NsCMY43t47P+tjKpWGIdoi3E/+xPkfN03PA6erS47WwNCrc0Ivqqp
NdOH69SDwkekqJAfahGRNgf0POKpsTx4ACb8xb1mSaglD7mZ32v1EI+LAE6YGyu6nFRCDMYR+Qk0
cHJ8iT7rL7mQcshfKL+bhcn575mGbOcUeWTI7RyAC8K5pAd9eZhzoBuSnhO3g7MamFfV1JcTw54e
6SgER8n9Y/Rmg9mRl99f+lWAukD+Q9CvXPRrXyN3TxYxXSKMql667jgcEG0NV9HbA3zwgDPMrIlS
freN2Fl8AV6UIcrByQzlZHhC+0i/a55BRm6fqFOnvusLgdbXpfvgYx06PJoM5w7NF3+JPwLSAPQv
EsLoD7cKB5EjmSzBnv9JNW11GNc2XprB8rtIu5Ug7jiN7iL3WSrEKn/P746Utoj/x+kHGlbsb1b/
+Dnm/hyUnhma5Mxy2b230YYrfksQzbo+wRFVUq6fnXd21BKZvT3o2ZC3SiRy3memUQypuAK7LeYI
Ebuh0NVV9a//Za68m+ZK1Y4s2BfK+aHHk+84y/Ekbi5oB+ATPqYYnGeIDQhObz9VIteCv7lcC9xW
AD4D4OcI40PzWZvbnyeZ/qKQLvDLc5au1vf2ZPuQQfX9lcGyJI2KJBmOEdo9tTWMaYiAUWfM8M+2
tHrpGtCU8uXAqIN5Q2OTPlCuszttVIcFaLfFFGsdz6j5cSiA1zvQFPyXm/pW7lfy/N/lcRUwOD4I
FhYdTs0WpQVffPNlAy89eTHmF13RRNMWY3ThdCCtjMv6sZcNc4GQb89ImSZrZLjVDCyCXuiQzkHx
mI00NjrY2Dqilm5orkjs4S/kjXgaNPd25NGmcIgFNkph3kjBkM1sMbQ5loCAkH1UtFwLkCQpxatu
oFH8FFUgwiLNNaWFgyPHaISaw+Vxs4Y5f9xXE8xwuH/go4zjJYGkjn37twJtlDXqoIC0RPeX+L5v
cZy+wbKK4gckRsB7Nq3P1gM17mdO2ht2YY49FVGMFj5FWtv9toAC8W7Y7882k97dnwQoQLQbDXcU
m9jAc0YdQFBLhvDW4B4O53zJU/CmLHS0Rb0nnRcGoGG8AAqRnLNNi/I6rusKSY1HH+hB5D9bVeXl
R9QupxRBIjIVrvXFgdb2FtXXd1jKGuZiZmdQN814lxDg5ICB73bmi7LdMryKPmAh9r7+Cw+/G+et
UymqGIzNmCoSY0RfKH/eh0i65gDXvxKldLD9siHxXrRmfsMIXsJIo7nyUD9vDBP+Ymfc03Zwymib
H6z2EEc15fuJHgflHpT0RDikWuE1GXBcSaLcmE8ykRDl6d6NlS9oViqyg4KUUUBuhZSaugQYTvzL
uiUXQ+3i0ZGXs2jVpjvh0ApL9SMhMgdRlOUU9jlrWATLRNB8nVtxqSTgMwmhsQD71GyeTdVIbBd6
noN2cTL75j4x+f2Rbf0EGmBRcHJOJA0/YoQp+F3QWDGS76JBAyTNB0r3F9SflHhX3fvDQM+UJpl7
PPC2BnkF2gxJYZDxn86PJkTTzUj2ZMmfA8f10250mqB45Rp/T+4lRQfJrcdcSD7KcLMBjhFkiYvA
V3ESdBTOLNIHseK4nCLPMGGzUyTG4BdIxzrodTlJli/mpNyFVXjEAl2akkfysN9EHw/3RavAy3ES
xm01MNuroAINitjM3PxSkezjfEpqwcojpTJvxBq0Rttr8BQELcKaBRXdUjDJC7vGtSvQ+sSixpno
JijDw/6KbkODfP1ZCJhkRw/qoFHKGKuB5chxtXdJrJvhGP1CUOMVfREb7N5DCsROIobno4zpEJ+S
CzCjm0H517gxEpNvG9lwJzdBEUFTnKs/bSF2N23nzYnT+nC6+NkpidKSaT7Oa9xeh/rDssNLaxzr
824fjrM7BKmEQ4y4jkJ773bKyA4Xermm2b7fGQviiL2SPEGMQwvtJ0AZGi7YQopNwbbdBLyeJuF4
vDf6M4q0FYI0HHn+dIuNWhSuqDiZUS3lPusPk2x5vmmv1hatTaRom54WimPVBmioIhZVVGnjGkjG
38GrGvvcHVF1UkULylUwpdlAX1Na7hrLxw39zgnvQ5u7A1NeEFT0XjDkbemF6ilojswVA0brS8dp
BUFHsSHlabTR9bcGlPX0chY2Yqn29rQVRsPDYExfLpDvaNl79DRj8DkX/TPuQwvKUmj03GhQTyQc
PB9V0tufK2MCJLrj7O5pKhbCpwBBZcoPtM/X7MfETSka6ygdrbbNZZSn8+sfMF2GfSrKK1yURD10
ygjCDaOQRbo8NwvoK8KD5ckI3SZ0ze0dIopaDKkOhnwflJqs5NIe4FJzsTAY3TOloGCpvGuS0XXa
MZEp5P+MFaBxYSTTi4d2Wx1NURvfDofNKzc/aZaQLiVx3l2lxpkZdONnVatLdL7VyHdwJKPmYjGR
Y12seO/hxLEcYmD/JBOfcz1276AJmr6l/ldBcFKJd1IX5/Lo8dRcFQrm+fM7VSJURwmtnVYSFoEo
ErmKsadw7qifi+w6MX8e0P+wQraEztCkSBx6siHCCMPUyF4RCWbFXTQoai05n0kmL3BJ9z4h3e8w
3WKaeOxtIQ7psd9oqg8fPxABGf+8pB4lSGEeI8CogP6eQ8Wb78O1m2KYJOjBcsIoy/5SjV8+tBf6
i0tK6pOGBDVR+oq4bVRbVuM+o0kDAcwAo2fWjUSX6Mao3UyPiJCmjXWB95t9PQU7x8qXMo4ndob2
NFc7u+Z59n7qeo6vGSgey0usk931J5/3u8KL38TCNgmxX5xLvAnO41f6FHUw8lDd5CLeIJcRlgQn
O7J0sibprMqr9P7m+Y7MtFSMeUnSJxZmuTc9lmktttYAn6DYgHbLinwcQsMf2v20fXDb2JmhJxIB
LMhchlxdawWeWc89lE3QDy7zign83a/m6QirKYJe2rZwm1Ey+vW41UPWSDdxSQhQVYiwqlFQh3e8
/+wJ8Y7Azd5ih/kPAh5b5EWptX42dSqKO80p9MFd3Ifu4JCGnJf8iAgbu9Rd05W5ILLWQhnonILQ
TMWL/fjDDWtV1kvgPpBIFYXLK5n6d/HnH4xIbTt6NN1uOat4V70243DSWdptPghfDqLjKKsZJf3t
DIVT9jakNRX3XdADUbgEAttHNMyCRBlFnpduPP7coIOj7FuKAu5QFgSrA6hZRgZTonwKEiMaN8O2
8JkwR7+CZe7pGS4FyoNwYVKJ9BuOfQPN4Oqtwh3NIf2lpr7mJrAVtUIJcT4uDz9v+3Yi3WUWm+0A
RWsMami1PowF9T+fB2jKG1bxSx1K95KI78/F17CT9CVNj0tb+uzOQviceMYYaYlp2jWKOWw6gWVs
0W/GHyUdj9Wc5V6csWBMNH1gZaGGAgczE43CdVoWjCtwx6zKDzU3o8tL5vUOy8IKMVSD2vkX+14/
xHipZRjRDC38YVPYTd+QARG3volWd8uSlxB/YeMLAKTymiPAsv5ZsAEmWCaGNHQKv261J8+pRC3G
1I+B2mEuf9TwrS097w2xpR9QsBwho9QruLkY34GKxoKEakQ1C99FSnNiukHIuxm42Ihf4AwkZz4s
xS5HgVD8ZqewyVBchdeXaY9Wwf5vjynEzOaXGYtz2S1V71Uqb/QOerZ+wgZHo6+9dT+xd0RrZ433
nak92dWGZKoeqjICDWeA49uM7BTvsfTiyNZBljAPa8PYsbbfA4jxdPYfcUr/s8ooTdAl6/uj74n5
nAyFJ3abq1ZISlhtT4erQURDTzE8b0GwQToOVdehrXbLf/u+sZqlNM2GRx36i+pOoXGaWzr1jxDo
hIEs2JNYh58rQPuI9gvA+eE9MnmsLNNz5/YRInvd9lAEIfrtDw9mHtVl2Y+q3/KmI/ni/bPbBQmG
9rt4iurNbVyszv5xLXJQwIYNifNChrdi9HvqiyNyS+yaLin5Sv0ggHWXm2cUcNVtFGRNGJ6oS5AW
dBNASqa9jbditY/04Y3Y3XV3IVsoT/KXQe5GwDIJ2HuEbYsA7bmVQ/ZZ2BASqAxifgIUf7HC7odb
uK7sx30cBTHbgN4RqY3zk1yhSo9tfe2RIhubMFRZqP1LCgx/h4BNbwOsLJD6iP5rP54ybkJ0LinY
ZWiuYn8i2+itXRlIcB/s1UzC0VDGdEl0PFkrrflMwigCwTY99V66Ny4WR+47DFwu0R8E2HU9rf+x
3Lb2DbU86duElcOCsszizdAoZm0Qrg3x5G7TWwntv36EzRHnj+SeaSIVJ1DJsQUV4NNf8XYEsIyW
qrVx9/G0g9jKJY2BWVFGP5O4uxIEJX6n3/9G7hnB+19eTOCcsX8JUax83KoQZzkesf652MnW1vnR
1c05rXvRcIWWD6lCpIyMYkyji2AgYkdSZjZ8oule2dQMauaMPYChwo/xlF2wEEKCJfIefjLRuDIG
qCwuoApNygvwnfCw1W/wHh2yqAYiUQ0asQWeYdO962rh00ezaLbnDOyJ/h6SgDdHpfF7u229m3G2
rLoXvfYQTTVOIdqlzm4r5fwDTr1FXrhbCMO+JvTBshBrGliWo1RjNSnZLk4HhcOnDNuLX8z+4Ga7
2JpyBPgMhcB1PsPD2QvxKn1zYigJ5YiKPVWdOqCeo8nADD4IeokuDS0sZaHjB67T0TFNQbcdCY+d
rQS1WzBFljuYDJON1BfwDfhU7429v3vQX7pf85LWr1Qrq1+HWKQ6t6RMXwgn3ehLpMyil5OQej/+
jNjrzvPHo4/ViKXWTUJgA0fsnNrcNxzr+ZxaDpCcLnj6ozWpulbivOOcAejQDqPjKWBcJKUH3MSC
NwHOUIs3JkWAg3F1F7bnqXA6KmuapueT0XSXYL7e3tEQkxIngC8mIOoynr/n4wPmJ7oMm4tYb00x
dMFe9ofXk4pMS8MRcAbeCo0I/A+iIrm/hsaJuTdO3Em0KXP9LzUE1oou5YavTbCEqVYFhMgSf1ag
vfgjXrGv4UuWgWB5hvySn3ZbnPix1XjlwbxSM228VeAd6VN+pn5HjjW0CXeXzQHP481w096VklGH
JKqAiJnhhOnIZ4wD2hZbbw28WoeBjf1F4LttiRpTdhhj8z8LNms76usfHdv6rgpMmqxtxnVaIMLx
1GMUw0QL2coZKjUNXBGhXKF2tBREYHVG9beAnFuQxZJtixOJaZOhn/4jvyZUQ2GSnBOigFFr92SE
ggNnLUYX+EdEFkb8uOnrQaqIJDf1T2n29/y/f6jSTKmSysZ9Znd3nOGyZK7WvDjO4rTHa1nA5hqJ
sTbD4ubDE+NZF/xk2BgTywCSMPSU2qM4AeEQonZ0DC5UhoKJNyNyEUZ5h6fEmwEvoesuhoCjIa3u
blVY714Esyg4dXg5sFaEjATyRsmMx4ne+DceQkfJ3a0lAFnDgSBKOndPXCKoe1Hu2xSi3ZFo6vc8
uvti53Pox0B3p4eLF4Gmt2B3mysLFSfOEguLu0yrQu26akxgxIXojz98GVdtgANRPHHhb+tYfS3f
QNwykQS/FXDFokGQrRS9d60TB2zNndIiNhhi1JMUl54RZdFtVaT2s6+j48BrpbRJo667dluyInaG
06NfwGHltPRLuNGK4XYxrbbvPbOLCUO7/yi/R5EIkqxNMAW5Q0g1YGXzZ7xB6nl24ieenqs/TXPY
Kfki04Far8Wtnvi/wudptz8S0CRZEm98AAMiRrUxTpYq+XLN/m68kNhadY0w1cUqCGJ8hku9l5Ct
28V2QKD7RW0qcd53O9KL0JezmGL0B1Qt5e2Mb5xiA1ZrPFIWxel+X6YmQTt7nFN/pY7X50CkYilz
oM2jZ+IRHhYP0lfb5ywVoiTDhz88KvWuqp8xZUIudSEaOBT0FVnuebWHumeBXZ9uD03cHa9vD3co
YV8iqUWfM0AfQGugxnBd/RY1IxijHBshv5K2nNUr+wJQozBVIw02Acicqv/QE6qnk9TtYRkjm0dL
zz1zaSpoCy0dPyKqn1Zvh78ie7/5Dm+/GWxI4KuK0FCPlYD0HYg7AK8Y1Ztvjvip4MXzmze78R8G
w7yYSPfAsoANFGEeI7KQPSVhh1kfSTml2/hxUy03H7S9Yag5BKetwUkGLOfPBvFPMr6JOjKntNFN
LjZO2nsvF0NxlAxhwx2aKRfCtbKLxtgxRZAN7bBwgyOSKdI7caiWlqu90Za5WgKGr9n3KyAb9TH0
7hCZEj/fXaMSxhtUrqkjNityNTehaTulgSLwnBMVVDR+fPUJZPJFE1P6W5RsWck99fo9vTZLanxj
hk0+hK5fku6cgqr3onvFXADbBTzhZgVvokAkVq4TyIV9h34SFlrfyj6WSYyhACD9jmM2Oc1z8zzI
4S7r63IOkOMx1Mhl5L5m8epx8vMZQb7kUM0TEbOfgUmaMrQr7a+usSVHN06XE8NL6UBpy5zsq/z8
Rl59ELOA/x6hmBplI3gDWObmdp7Iz63rGGgiyDYRw82jN/7g8KyEiHD4bjpPBbG6/dQ+Q1crTYr2
iqrVGXJ6bqCKA5iy7C+0y/TPy74EZh2rUpnUjObX16Gwtgh1FzHJxKqIB7LsJ1Yj40Hd93QXjZK0
H2Wabn6fdovOjMl28kaUS7aYPPpN0cd2M5Yp/c8x3St9OrJhvYuSqDByCXBiPKsMiznMnj+bvrYR
+OKoKaZ2AoJNAL+WEg43YjfSin8ODVAFwPUIQR+L0xFx8FND0ZbFjffS3TA6/lvAhjznKr9uzTyV
pVKjzH299BhB4xuCeIMp009Fuow8z1XirpTMpgjz001jnrK8mtzNZ/3QefAs0KgjbVCO+6iyYduw
CwlB6vkdQ7jGnV0lnGFi3H9I34DkuOISrx7zgJbXsrrKNkYQBmiYr3iVASlkUwT2woMh/vjVCco0
0UI0NuRBwB4s8y2jfSOYmuz+V9VJ84ozRDByiQIx8kbtMX7OOBt3+fHfUT3rEbI5lj1LeZmDMutX
aydHqtWfSqkRm/L00+UARW7kurYuXfQvraDIF7GGDtnWsU5t+TZSCSQsAIdDgdM1ggK0i0rE+5FL
rgASO2WDDFWhfOHI9uhDosy0Ihh0dXF47IOTnVIPTj95LyGxlEck5cMHUOIElIGnKC8x93Jdn2Ro
FJTXFe7c/2JuMROzhb/7hC/pRvKXqdEmbJHtb9sJC910Yw/URgP2yhprqCzCw8qFiogMyEOyx+00
PyJZgk2LjTHJvAA1L11K8BvND49ySFI5lk8km3YEl4oGtwkIScwdIDbcEhc0k/eJY+LbBIH1LImc
r9sCfkiov+y8bVM/azHpUAneL/9He2258xwnpT2UAEWjWBL5HbKfrteK1hiIa/l0eBOcaMsF2GV9
MZQZ6w9v0biPruQ10BR2MrUw8aTO09IfurooEuKLTYXSpidVjzXyhRHQ7PAzBGAShk60MqO0UoJo
S8VJQ87U7k6lPsv3gmu8bULLeaf4e6ERkft2Lxl2qJFZluTcdMiLAjTI3Vu98/rrOvKwJS3YIOdK
C3SiDPGtAI1QfQAJASzg7YVU2w9Dm177TMTXV/SDgIqBRrkQZ/4N3ClGPt9ms0hDSQfrs2FTtVf1
Sr9IBthbVgJHm4TgbZXZ2vUT1fPMKIr8Z72NlH4OzmB1pM/XRKqHjc8F0IqPREPF2bWvy+Qq3lrK
n4K4CT9o20QAjhalzoejpJHor7m9HEbXv8JmTyJVGDnlJlhm+FoTSIroQAi1UNSlQb+4vMnSkfvU
pOYJCq1Jpj5KO3ZX/CzZnwmBfjzYrkCBFodGbzj4sQeZwfG8sEu4QgtMW2nFTBEa1yTa4xnjwbJr
aSoSvuqIBvuwotrpscvY/4DXe1gZiTlzvIWbocyFvV1tVXxBORXAh1p+HFLnxfHaEQQadjDd2fFD
YgNHdvqVUhLlpOZcScqJ4QKTeckMDJNWgwLPcOxFWXlHXsxbk6Np0o9gDoWH3t2tzaIPONmdu0CK
g6EBK4NmX0qPRaZ+jKCEpOB0d3t/E+Fa47gJPhyUNeYqG4+3Lv7AgYsYG3x99WnsDLL1LYjrgI91
lPtWN+rErwhCPLhHjBFbMWM5c9vnhD8BIaH5bMgiDb7wNT2kMIGsccismAHnQYxFsBDNO0p6FHZ1
SG3QBZ86/5qtGxX/nUZstrCev2YVg2AJt3ytEe7YXQZesXItEfuj+wfZHPzdGwJ8JMAXd6LPAR34
gKyUpJHJIzPD5o4kRW5orfHoHi2lDqywtenzTktcao58dPW9Wsnx6NQ6T+Ltc9RDAyV66WytUsJG
Xj+CIdrFes2VUjhToug7aFpMg443kF/K3iSwbh2ErU/ltWkUV8bNku8fRjNfrib/hXTPzT/4tcM8
uuevG1Es7E5lFsQ0jae5YFujMRuuM3kp2uExIgAaShe3TnCA/g8rw+I6JPnN3AJQVHiqh6ceDrV9
zOPqhmaiLSkz4JEZvydS5WwpyFMQYBRNiVJRdieHGx2TFRIN3FcNC9OmIzvIiO8fYwVgm4g8jiv3
4HaB/vhSHpNI8vUYf8GUOGEyvWf6XJqSuu+tVflLLneTDo8a6W8MrcPc/fRpWxfYIaarT4h/rKZT
RZ5amc1SyKCArw7xK2eE0kZDP5279HhvEmyKa2YfQIc0KNY+4y5Ts26tJiuaCD6Y2G7OYWHnBcBv
yomBW0TVIcaSapdS3UacLTxqZFj5uRoTVV9G4N+mICcKS7ZAZX0jMkU7RJnfal/bBT3XbXtyJPUF
BA4s9rT6x580hJJOYutvDwHwxc+XyLOF2opwbPefxvgMAJ/DJZmw93Lmom36LWwQ4EFUWNX67xXZ
EgC5sx5y2dYyItdv1DiTBnWWU+eT3HG8y+D2l89O4JkR7pKDDDMZYqhda0obmWtURWaCM1ou27n2
CQfjs0nV4DWv7uhqB/bI0Xb9/zznUUhhCb2WIx5aH3mgr5e+0vAmuAVOGxguGlz+satdL/pbczAP
onD95DGxRBmgLdXPjqVBOwtj0Hq2mfDOpNH1Jaxb1ZA9PKmQbmXDnOk+qFoPYj/J0eH389ih3ydr
HSFS0KRoTdylmcxP40vnKJFBQ9bYoJ5xLnWbzhnkmGX/67rTB7THqunEp08uRnqCHM8KzMvXx33p
EDl5nOxtgTE73I897AXmUVhzaKKOpFcH2w3eyN91zsY7pGp/khXO2emiiKw7klSHDyB4YA+Rarpr
+ovnRcl78wd1QgxObHj2VaWRTxZcLR3a+LfWj3WcinVuGB+uHCuKRQ9daAeOAYwx67Uk9awyf8n1
ARZjPYE5w7bveITYO3W1iMmzwR7AmWh4UdT6tEFC3b89p7Z3ovGaAOKB7YJuoL6Er82zOQmSt2l9
UVc6HR0G6+LJtYep1p3UJP0OV8XaXifElyBrTgo1vcrJEYvKOmgeUAWderYvwyReFHK2+TzJ8Il1
N+GH8rbD9e73ry4lRKVmiqC8wGgajyiQqqpXpnQShLLv7rc+TOHvENFCdX5aQOzn+6p5dUoYnem0
qJvc0HRgbGPmtzpVjtzD6j70mqoAe/9jAyB6AVxeg9kdOEu/VxQEjkuAYDvk9VyF+cSvByGFyfiH
9ag1hkQLyqhcpIa17TEPp5hbsIcnBSEVlNx43wmPnn8mKO73xO0OIyEMgwxx0syatAjENZ+P1DBk
Llp/aPtKEqdqEMezg3oU8RJ5f8G5ygNFa80P0qvEYUYpfuxvYyAEYB/9Vz0GL0w/AuO56c3cnL8+
6rSLb0ciy6o62Y0JOZ3hUa4WyIbqdWYRpWRi9EKatNXPz7e0/9PfO0MQZRLL8c62nwYsGqJs6C1C
UpqFFVDQIyPsUdyjNYlA9QPCxnPDQReZCeiZen5QZ9mViFN7oxTlhNxXIemCGKJr6ERW5yWOHrUr
cZGcyhoN2pd7gMDxsUidX3GFokdjncxnDLjM86EDeLjow/HLKS+oYkgP+bTGPxa2T6g6u+9Dfe0F
NrS4IVz9o52Xh2yrumtm+TMX/TCYk/yeoZ0ywN8cGU1alHTylB1XJvJc4g9yAAyJ9QQ6+Okj+4i2
y3TEdcP6wPVloYeuJ6rM0JZojQnkkFoJh4jURbWZh6dhE/LfJBdoldBiaLnVSZ5fBLpBYBWC+4Wv
bCchoFQ/m7oNsb7E08ioQUF962gie5J2rXUJnQzQJXk8M2XyUI9f+8Cm/rZA0rx6XbDrdSG3suG2
OwbZOeB1ZSYp/Tgq4zkXqfczd9zHBHSqhB7/cy+jfZmgzxmq/9YWgaPDFw2NuG4bosqOu4RSCa62
KnnU6voF2PX2IC+eqJJIydN3RHQ0RbhCQ9okzba+VmiOUge8vvQWvkeFybNSP4FFOQXQCLSu31Fe
PniHN2WMw2fxegl6GfjB33Sxr0nzy6YaPQT+iaZnB0H6LqauGvsQBLBXAKyZu5nRP1u107NZSQBD
Ru3tq7zmgPHP45037L5jTxiT/T6i2nDUZX7K/j1/FjOO1Yy6HYunWQdznQM8pUAHXmArRCzWSEd3
Vz96dUjn7MSoNwhgR6KXaudyBXZAyIabL/hrorQRz0PMEsPigO5LCVWuD5wN4tOLyCZ8dW55oxn2
rgelIX6Xquv9feUrevH8dx8L5Vwkh6dVhLWTmk2C8VBTrlUuFtVAS94fydcHBddl0EDCtSg0nUkC
GDtCa76ORoU6vrL8ul0Dqonkxl1BTetkceKV0f5bm2BXoHQCETZHvqPdxE03YSvytZVPkBKZhuE7
Ux5mkJhEUHjkv0Q9918H7nCHWtR6etppBsfnJ1GjXHgctHH3OemXXhX/2KaQUM+7ccaNwxj5XB1P
uXtMh3Fwuoi1rYFk+eRT05kLjlbwEJByyJPe8tpmmIioCUS0wDXrffXNesbxSgzVUB2KhPVPi7hT
diRaFZ/jCnr6LUoTE2BqGgXkusLHr3wbbCpDZrYKGhisLwdegdSDluvUtD+ABHf6WP2pWd08snvh
3hZAXNjimTiom4qLyEPtuLk9CkPcNZ+pIG9fr8je3pfhDZDzTFJfzivrT5N8WVReYWAZ5WdNMmRo
b67Uv1u1yHBQv0Ea+iVh+/yWOMwVFLPfT2F1IYvN5lQQEIiuG01aYSzJvl3tjiDYwPp0RribndSx
yStR6duz87Eyg6jq/61OzeZj1zrSMpd6ey+bNjRf6oq1Sqc1HPXE7MGmoINJY/ZA5bQnuMzb+1Lg
SvSFtVuU+6t6xpc3XNFxiXHfxqiYfOvash7lUoyRF6sHET0NL1rjT5FDf0sS+56KMGts0FXAr6vw
BazFQGOYbjpjS/Bm1vZKP1789JtWlMMU8XRDi4E9kDHWQZYy2VJpgb/mY03D6GJfjeNwOV2Z52W5
RSyDGo8qPfJz+O8sHH71uyt1YsO8DWdMVhoEK0hCNnQpC4obkI012+bfg6tRbhK7K994HxnKt8ti
v6F/wNFMMudOiJm7K1eBKpERrDNfhDVlOBUmGLKGtjY40dWil2BSl52pD/wk5dm2lw0LSB9XLFyS
kRD1xV9tA6++lDqiTjdVdq21rciHGd23ie9GeRFKT9a/MvwTnPXcgfVOJ5IrWnGj4Mz6mldxsent
T9B7xJ+mV+1zlKLuI9xwbetptsfVIyntDZ7b3sg0igQbegDPC3+TMfwW5nvHZWYweVyeg8Pwidc0
0GSAc03UpS3UiXH4S3r2GXJsz4dJoyYvvua4STGcDAyag0KXzCPnMyzQzMRgtSZMPK+lEgGz9C0Z
VaCo1654hObKDgbjOPuaaY/cgYyOealvn9HR7hDLgMFHpKC25YNmnPAXLnGS8TatUuV/j1Wzj+A6
cyhKccbBIxBfhVHFJGomzQi/UGdS7mZ4iBpp2T6UCU2WHpHyzYG0pY29LUCqDlph6BUmwnBDaTuu
W91MWJz+wpWODfuyvISi2+T8lni63g1QJiZSuKHcWTwt7AvbmbpPVgt647Cdo5YV1y3Pifk0wJS+
zFEPH5GkhMCKp6UAm4CHbI5jBZPqmSYiNGO7oAIzBRq3jTexhNiS8THg58/u8IuNQRFuuivJ7uYo
vvYO8Rv2D6TaGN+JjzEiuoOovmEkfBPiBU3O5s68irRH+HuB0lNVdnWdj0YH9ROWit7Dh4zcRgO1
JiYWhs1nMl73cl7qeSOMNQRPdesYpSiDO+A/J1sPuRnTnG5CtBnRue3wLXFOpPcHVQZZ9L3+sVcN
oM8U/KWwwJmUBTCnsjuFv08Ty39uGJ3ttergbUB2aTYosxSkjwWkw8q5O8M2OYisIXO+matUUmpp
HfY42Jq2Iyssco6neqOAcz85qMS8WF/BdEO74opAZBx3MGvVra3GjQNTtNlrcz2RvGhby9tQhcfq
as2mHJoaZ+hLPF38VZ2xiOHKLt4I3tVuHYWIF9TeID2H3JHrg7b7rrqz/Qmkp+yKz0grlVMp3ZGU
gRF/vIkMjiEn0gb97qcFiSSJtJsuWt0pLLFjTiqXm6NaQpiQPR0ylayuQ2cJ7tuh6HuRT9wLxKGj
7bleOCdy69cK99cy5bVrm7D9sK9PozX1EC4CibpXZ9x8u1Z88/O2pI7EpsSy6JqglcqKNJGIe5SI
mHVeZWgthvYcnbkCyuYh0kZ54AZi2yINbq2xmcRs9h88h7JiLftUZf3ORph+4LtOYwQY/2aQLU3v
WfMouWPNU3EkgesmdhVIW3cRr2BsSVol9HBiGVHSli3RHAqJEy2WPmB++1hWNLNf2/x3TEgSR+8e
Dsg7tTRcJGMdnt7DWqqju7f74DFpAy6QCKv8OjBUHQ71difyUojEAwu5aP9A5jRKiXYhU/kA4e8g
oRnwlfkTHu8hO3cBw60DlJ+66xvNcdLCDRC2IJvRaJ8yyQq1dhzAc2K06y54b1tuh9yNxdU6LA/q
In+e50HlvABrq3XaWLkgnOHYCEpXuIJpH3LNLKkWLLAypLj37fJTjL6T1oIUOT8CDP8Nca2VA0Rk
120Y3k3LCVdrGuBlUWcRwB97TcLoCFIJXdxDB9UpaJmUENjj8Z7X2kojUbL+aJ3dMejkSWyKF6S7
/r+r19Y9is26xDblvNxm/bZtH1bg/KgswR8r/KQAaRzlFd7OsmaytGuRGShQ6OMcQ+oKWoSdk7EN
KA06lk7Wfr10MhwsuGzsvRfxQlULIMxzeoFfAmpYVnRrEbzNOnk8o/GV9dKuTOIlsFfn3Va8WWiX
jTUAJThsJ5J+xXbGiD15xbxt1yWE3gNVJTr89Un9tI9eAxB74Xg8Y5DMHz8wr1+i/4mKP0yCapRs
Mb8+ezhkHTKEBUwFsT4gWKKgBVTiUY0SkyuLnBlDIHog+ehQRiabHYSY/dJYNYq9aizxCCMOtHNp
cmuMoEnt0eeOxm0X4ohlulPWMMvN7LnKwmKQMJh3Pyq8VdDBri933iAVuTX/+pdpef7wRElt1Nlt
MAkpHLZ5hT0ECChD3+Dis+U3aT0PJfVXRaMuVWQK24Y7LDSZEl8rs2Reu85iFcV1XsLpu82Wk+Xy
XNSdEdJemu9LGhr1yeUSwfhI0YHXagR5r7dx2wIZO6qVU/IG+9rQvy+g52GzSUAQUCjiIK1R4PcA
hQSn8dOu/qLiVJG7KXD6UJo5NOE+cOzyufzRh6b3CPk7x2FEEJt/ls0ej7nYbFWiMjACUNJjUpsn
3/tcIATQzfmKOp/L20qS2W+5H4J7wKk6SnAg1XzYCdHgXMIDNJf3mrr0SkpOHC/4UbFXCvUxSwkB
k3MfAV8m/P0u+fD62eogsuixmQJ/OHY5CW56UoFYipHsr2duo7NWphc049caqFNtuh9IBVy7qVL0
wTk1K/tv+nc7s/DAW6xwEXkwcldV7Tnx/zhOFFY21uJVLbXr+BTKAX8yBRHGG+DMmCpW1mS1NNlE
IWARwpoV4G1knSwrTa5KbC2W+NkUlCdsbRueVaHtxB0gZwdC0lApIfGkVQ6iOypTVZdwWDcFrUAe
kHGD8TOj/nzJ/XLi7JluZ1pyFUNtj9UQmW2xyjPSyFaMv+zVTGpddu11kYGStXx80pNrOnLwamRH
NOl20sct6zSjr3JhETDyN/+pJRJcdM3Xvqg2cc9EvTlq8ncEuVJCy46bPndt4DcA7fyIutczjlw6
BLhnGd01aL0da1Ay0a7KtJCm+r4gkP7jxCVfZzsO0T5c6ANbY64+ywmTO/SHwJUGLemuDoK74xCD
VRHeyziXsaGS/0NfaQEAfkHHqyyA8NHhrfur51Z9wKZxVAo3ouZl0iSwpaLpkq/Rx9IKPeziLqFk
Umh79KgaSoH0FlAS69Pfc5V+qRAxWJ7yr6NGOoCNv8O15oX4FQzksy2FptWQrYVkj3MsluAnf/oJ
Ce0boAIgZA2xkSozCr7Hs6xdIpX2H2m4hz/UjR6gVgDaMKPXTME5oncTuUysw+6NUE1KKwaq9VFR
/JKczO4QwlkdQD7jjKBnSG5ljfvNU6ePGQR4SquyDWSL4YsvnFPoVjQVUwtH5v35v6j9/H/nZLEJ
lhDJ4q4pJ3sGL9oc3KEN+eck+ulp2On5cNffHQEp6r8Hz2SO6N5BeZIr91jYWFEjisTjhsoxWAAh
bxnStsnoLeKScERfdwLiAhJ8nMjaILa7aE5dIc1TMyk39+Cg3yA8tUySTS8UraNdjVqemQfmXWAZ
vyHxaKo5O2I7myXb+UeQnKhHAKDMa38UP4q8kCNz2SIDBfSQ7iNOEScf73aPbpiZHVl5jQtA3FCr
tKq1BGeSSP8trM6WHZmzNnkbXjdPw0rjmdUWyvNblct+2XlfSSvCF8Oukmyuvd2gRed65wkQisZ+
xeo55ODd7Nv1fCYMiWEyx0lsARv9+kJBN1f+eCiIurJz+DNbKFfIKMzy0rxmOy+4GE9kXLncURz8
IhE1q8v5zwO7t44kqItr2oHQnYpo5bnEjvOgoP6y5ScrYLrU4R69wpjh5X3+H2qNCHl0+lTlDhQH
Vqczdpjb6U6BMpweEJI5mUui0H28hcfeYb2BYcCMOb/27tmrFmz7gZXQ1FOfjgR5Y5KE/FXJZnzi
p8CqTTaWcIC3aivUVQ/NA6u5wAWWnkjUfPfJtH70wPaGcom0S+xCTkiyRdu8WxMLptZF8xKqEHpS
oidbJVV4EMnx+XufoJGQb+MMLClkam7bhYB8tPoUmnLIxHd2KWPfq7N0FkfTNBjsMTc9vV6stsSC
xGUuUUBTsygd0SG9gZnoJVcahJ9qW9O5+yz7o3MLG3VTmXUG2AFyybopbWcBQ1UHNdI2FRjNF8Rf
zsHC8sPzexMIpxf9JGTXawHciq21rvCopdUQbEXf4gPTcfUhGknKhhOFv9y5Jy0mZyBG+i1QggiI
Uqp1F59X/Ifr+Cxjwqw3U22dg40azbYcuYOGjDAy4LqmVrAAky5xnfKjP8QfUiOKnpeU/+6wsTEL
AUjp9pdXTGWM7m2r5dv2KA1UVNbVjQAJOQUU4aseNgHutR6yOEOToqHVO45EsiuS49Ave7Ci9k2f
zz2xTJdjThAmsOalR7b0n+vuMO/7AH1zcjvIuQX98jlCeV67rKSUWFGgQVhrLNfcI7W5gtpwlzUi
Gd7Kvtut7uazKYsaZ+gI19BdrIMHxiDVa2f2gjKyLUjL2Rwd+Pvn9O8Bdtm4b6BEKb9OFzGE9VrQ
OwoXVp8pYnVJ/B226Js2HNBdJLKa+wT4tm9mKJB6+yyvgE/7ksotVnFGosIIcVfqUK3iigtuVaGT
99Xd3D3VKvIJTYTIhy4MUhB+moEopETDp/Ug0cwPIjSCmgHUbZIXHcdQViIL8EWP1cRVYB1KbWV2
XZ3QbJr8kKzphAZeVM3s2NP9E8AnZ4L1zFiOI9LVPXVl4peS4nFcfrmIO+g84JPgeYqTvqXlgaPN
+D9J2oGQfoBUyS7dJvh+qtrHRwRh6SuT3evmlIWxPU9u3tOpzD2SIp9zbo/nU9bVE5zpslXbAiBl
/dOmIOpT5vLbPhVNaJSIzHev2wO+MGL+M8yGI90eMTWurMpQrDPTTxI/pS+Z71IDBjtU67B0zfFt
HZrgPhHzuJMCQhRrJxUoCSFBLfd9cDvnZSvnVyQOh3hm5S2iUEE9dMBjtbpTuO6nDTQWmj7ybYWC
ZnaVVmhN99HpmHWO56h2i/XYZAPjOpGCUOsEXZdUmKyW/PEPB/fX3FId+F0d+LpKG+mcIAwsJv5Y
j3oYvfNqIdHb3YA4zjJzu5bZs5MxuHsAsJXsNREbcZwDa6llF0yOInDyirlK5nYAGDXckRJqy9V/
8vxe8nnFBV8eblhs3v5xm8jnCo/aTguvd3D76NCRnkcR5V9rxAHwfrAgd30708xx1ZiMjl2Tj5Zc
McwN1SE8M9vrgLcubkpFmIMX44lmXKQ+1Z3lBQjTB8Aw/+hzixO97TLeT02dhvHMLi47B7zPejEW
GpktoOpWXOgET6FzlLR4nwheWVqrip+TxKyL3jeflBj1iPMitr9ERhD1tdGqw9KkC3SSFB5Acw8s
5IYYxrQrPCHW+KUCOB0+KMy90VxKZRizJujgpYkasITTPV1bfJQmPqwsRnaoVFyHVDpphztOmcST
SZmkrOydkr0nhhGCmXp2lXuVTe0c8p8uer/RsdFhZFb/pCSomKS+klpCgedg/7GUIYqv+j0s4kFF
jJ3KRFUsTqFKvqm2SKUZgKSfiEoHB57yYmI43Rz4oGFPTKiNR9hcDOdujSKkbhZFBckMde+ZO+Dl
AVsQpvJ9eb64g80POJHvtOlqI+OcXJNkSaKHnS/2ABWZ5z6g0dAqcnrW5oNgGKpDS1qh5xxEiMMI
B6Z8Uw6J/3vNp+svFhQvrevjMpnOOIYJCP1YaQpoygSLyVspdBNHC+pKEixLPOFu0kjYxBy2oFqb
PeBFmrxXerKL0vW2bfaWTQn4PDQhWS+g6ZeoryHS1GqSf5LkXPzVTFJ13qyMXtpwshN5Lh5OXus7
YUHkAFC6Du77NN85CHbrK5rfH6GEzeavBhc6jxlHTq5fwSldbGADiy5G9byueJSG2hvlXPNatAzB
lHICXNgoqsSwtcVCBMiPJx1PfnWgybF+V0/hgSXHUrltGqQCgreBMfaUgL0dmr7yAN03NBiJvjK7
6+lXJGHq6vaeUA3ySzHcrbFPIYoDlrsTaXd41hJYzImKmpVpYQbAg4WNtHjt0FZ2+Tj9o5YBsofS
TU9Aw33P/6NBL+ZTN/9dlldCMLuc00TV8hhwJM0Ccpmg6q9yY7Y7Ov6/JSPbAUdlFaIcZ/v44Sfp
ecUYL56vkq0uNYM/hb8IEyBrJ37t6E8OeYYFJiogRkmFeFw2L6JEAVjifTD6G29CqUHjgBJMshcd
U3h9f3hmiuzI2DmDVII5t2flt+suXvHFcyqsl9Y6H00HQ6/rcgNXf2LvyW8P4lphqJsBkH59ywXP
8notnqaBdupXXeK1uGedSBJlPBSc47PpmR8xIS0tHcwS2qZ4rT2SFQJFNmYR4A1c6wq1VPRvuXCY
KqVdp7CFp6nsoWMpFr2SXQzVpbmq51l6THkpDE3TBFT21WpsPFV5t9TeobI8onFUJO67QbUqaght
e062wTwgdrPhsNdV3TsEqnM2JTt/k31aQN3X6aT6iwGHoS8c3H4yNcblKQl6mSNXnxITFmsYU5W7
MjWIMsYCCVkuj9EKGRj45k7+GTcxYf8NHEuZutrTs68nipT/eU5w6tiQ8xHz35+GclzDhgyi95zI
EEIgHdwWVUzBwzfa+m4siLOGw07SIIKx0AoS3PhVEC3QMXo18+1DrJNDvIiqoaJL5MWjsl26oxTp
MKZ9e1l7Y+dUSD+N/mcy4YEXsVS7LRCjFyHTs+vM5yrlWKNQqGsG/L8XGvXO/UgsRB5i7P4akQ7Z
rWW3MbTCpfCbc0usLYDb1fijPSUBgQ4XlAvIRCEWSY7VCPkZWKsA3NaNWPoZ3zC30mu0YWxpxa+q
Kh9zVoJ12HPiMsC2NAH/PthfVjxqMpvby09gHVt0PSgDlqqShzDhaPxofa6zaR5CkC6iVfe5fhD2
/U26nCCuxLsD4cnKskYADnBMp0IRtjvzmdusig14xw/tM7cC/TM37c8kZNnJJXaTXjc89ol9CZzi
yyYfOOb+rVGhUZpTok9UgYvtTe6nqFmrnuWImRhJ1PTHmUChkamUpZexjASR297bl/8IZspV9XZu
RqpWvU59VUeCC9BBiZn5PfVqi+rBG6/fKEq2fEa4f5DER+V0CTrRjlN5uLgXTmjAAayFgfbqmBk2
GEauqTWkd4+JzOCevur0LIGuUM97959fNWmLVxS4AVRRxsRveHZpdQV0qPsWh9Ycdo984xLtUbtL
Na4hzztTRvQ5cvHUmuoUE1IR3sMBO93S14PJnP903rClILh6UkPnBBywoYKRDo+0DbKL6L1B2I7z
jcQkIBjFYVFUxFis7pbJUYbJBR0Q0Ml3HnoOH2R4ZxQalZe9EhnpXSj6PbskRNBFlFvYkv0s69d6
becGQUcEKRrStBi5Ie3Kyls1m2755Ie/MUbxK82dVhURDbyEKYN2bejbJzN7sxxkO8bCgAtNjC/y
8KtGPY+I0xSUxRYykWC31L7p/DqtMg469OO0iyXGOS9/RWxeoeVjwHNWYJX8erqUmi7oImbwlrAa
2qiGxXRGWN1W6wfqeD1D7FaLGlw8+O1P9MpaN44Oic9RkFespQXWiZIuScBp6M5jPeE+HY/sZWlW
rtCUqeLszCKm/ESmxK2/HvvnXy+iXccR80Gwi8Fv8cInuex5OI1klaiD8wfuErGXP4QT2B3saiiH
4O0gsjJ86y5a82zotLd2iVgQ37ODNCyAKeG425f9/FPju3kS/BBOp5njPFKC9Fr7li8I6t5TFFGs
r+YYew0oxO71XUM77+NpgB+gwJwSXms1dl+aBZWkFU+cKztztvkWMIqfJSAJ9PCLw0HlvJI5fsiY
GTR/sWGIBiNUib5aTsSpx7rKGg1qQ2uhFkxUjeqHxC8bxMUC3epTyLZ9vO8jm+2MsJqtEHqLOJaf
oYxfeE3v82XOdZWISoKyL7pyiWsWtEnHWRkJMtpaIZkW1dvqX8mALn/dZ7anNtI2BtfSYDfbRDJo
7/wHTVODnZvygcZ7Q+DR/r3mKIhgxnbnqZsX7GXoVBwcZnTMQuSGLfGCZq+vnuroYztuiGqCda0e
d8ep/l684QWpzdrWsBrY9MQGBWGOZuKEnwz63VvKaUmT8+2gVrDsXshcyfxTw895V0L3N5M14GjI
Fy/dRMgeWTo5sS90Q/6zRQF0Gux2H/rpoTTvoTEgQyhr+hKBCuLzJycpiDvwRAyI7xPSLIQNS5fc
X8z4HxcHwxDWrNgtFZQe08AZ2GwjXZqiXlCtsJZli2cTF4meeSpstXda5EK1NuTZvxsDkneRHydu
aL9Q1ssP+c5MG45Ceeoqv4nl26/a4PaaTFbNeIYiG+Ueq7fu4QM5EUW5Gn4db9Fjua/tKKynytIf
z6KoOD1DQ+DZ4/AoCmc+EyldPVFcwCBmKiVPQqcF6nwf3k/f+CnkqYLYw8dr6j6qJygczHv3WcDz
Wq/2EmgBLoi+3Jgr2O3Nqv6ti8nrLuBn7EBB7+rrbC2/8M7DVHhcN4/Wu+p88siB3rrpObMjOeFL
Vbhb1lJat12KB2K2PuJJ4aVZt+Pfh2VvuTK3s8tylgby30E3AmvdGYLATVmoAfXX7sFU1WwWaUx3
RqhVZn6TrPDxkJeh0NtSyhTQkIwjMe9eFfSpM8+OmQdQu1ib1LUUPxT94fLCczVPnaJT/7zq6vlN
evlWnAmVMUCc4PmvaaEOcZrmFSe++wm2k4WqwwxHzac7apur2tV/dBmZTuzMS6TI0vfM8Ld1VPjK
AKNXCDpSDncO/4oxdQ6HnXdCHwH6CQFmIcJQp0XxmGHFWJIQ2lgrlTnoPrBX0XFNW6jRkpoh97Jg
WJSUmOG0ysRKyK4Rx+aJWLx1pl4172pJoGDNUWRiiddW9fsOhjKtEnUVak3XVchZFw7AADQOyXWQ
3/5k6nPyjl3fnnZQR9kOrFrdMzmwSnN6TqajLywlKephO6TU7qoStCuw0R7KONQ/N4JsHIiCVgvR
31UpwtGxZCyl0AehdmlL6L3HQ671S2fZbm0RfGhg1JFwO1riJ59CBqo1l2QgzrmWKMyulb/ErhzN
8lp6okwftbGR2JcAvteFhNPU/1MxAWzZOUiYq88x8WOMMwLkefgDrvxNnc719fItYXZ+CmWB0nsi
BPgTnoXDCpw3q+hAZPzFwIVy7cCOVcZh/eNKTuGujIHWBgeI1jWwRMEsevz/qto21Ph2ZBKrt8FO
+m6A38rNYkomG/QpBK2EfzFMB4IsZ+enqv3hG426Cx1LinVm6mwVV6Xe5xDeuHx2OzgceJBl6+JZ
1ZxkQeGL1i3/jgigxQgjRXWVRg3CrF3wt9kCH5Gl+3gXKh3yJqAxZp1310bLWN8ImfXA6tQ7CC56
kf+US90z9DOLXw1sv+og/xuu8FecHaKVua9lUqUSpmHOuS5Ccm11ZI4gcGya3fqgF/w2gtzkvCVs
JG+BWsQa4eiNWDMxjOSQex5ja/0n1tR8ibfz7HBAWNZEhHV7mmXs0gpXlRB6fWiseSEDYzs3pURO
d53a7/1tIyrLuSpDdgwtwOJ83rgse3o+Aqo6DscxVmODHXGBBCCE1fqfeY1l2fbj5CC9dmKMutc/
pTfM5aKE3oCOHhLYyXiwWeTNyZyp+vJUUHfowcHtRCcxQxZ6/cGqbL0STOIZYpNTA0+sWornZd+W
bRhLR7QYbPPscuouWdDDkM8iSlNl1uGXzJWE2QIxMmRH6IHbEXkldM/ZejZ0UGHVGJQyj2DFKj9C
pX5qdHnJE3GXSGLpzmKhMVt1apEjlWU+nOlFEoIZ4GKINGvdQq7jElammALKlyhoCctqgpso4YWv
VBhueQOplXFwziGykFQpdI3GUYoA1vzdA7kyUS3KVKy82BKOTKdyE4mkh7r0Ec1TBdaxIzfmV7tF
dmkNmKdH+RL70rZLT4aK8So2CnnGkHj6iWKN0noTDOvlqdGlgn3ijV32OHM7glBIj/oWfFHFMc3K
rLrF9zGyJS4qsPooiKxZVYMuItkrZs+dK7Tk8qlUgXt62hOPQEQVFyQbTIJzicPdMkR1t1/fUhbm
hgszjmeOvepCPE643iRCZLJ2VV428M/Nn7F5SCz96umheeOsUg4TppnoncwszqCMP1dwykO7hnw3
VpITGJ/iWofitiGG5XEHdNFB3F6mpGeVn+rSMeLhdnTwBtUDv/gFAciBNhiK5OdTaqdX0gPDBZSV
MGjrzbamxkfyVStoI/L1P/p9IoeM2iICMAAPyuPvXyofBC/ka/OePYeALPKo1wmTKkRx5ywO5PR4
hw/D43hLeI2hbnwacyZveIqq1ksVXkyoV0WX9HHdA/iJDNTgmc2AhZoyO+UQzb6jSQ1hSo3hTyG3
essar/TJnALagqz4ogr0hQoJNBED+pNIH9BkD1wzxwJGmAibJLXqtnjFrzQB4L9HEwfxkR+RyWYf
WOT3bhyVAK/a1S1CfFTzU+TNmPBCHQPZVPUktGsEWTv8MBCSrATVfjeRjEp4FHmYg41oMTA1nC7B
B93OHu81xBE15p7R+bBuFzeXALRE6mePjywNR9ISSvVDXQo5ajlznAo8RGQGCTNYNAKUKNLuYnmz
zAddngRcJHA8rCk7iDaq0ZwjadAfJUm2JlcT9OIPTVyKr+We16HwRN1p1E3z9WqbQytQSzUY2gHo
wurOnAi9/OBTavBdKBK5sDdQTCt2M+DhXzZ0lAPPhogfTbwnRK9o33gjmDqg/AwTjQKA6BP5Yasy
kZYAJaNXmnMBYp8OzF7iUfOYIFhgM+Wt1Ujqr4oXoNjpI1TR4yJjZXiY55fhRaopyMzWp2EHzzHy
G86IzENXAKL6zgplHnDYjNAYyWkeGSOVne1a7YbkRh8bBPgwx6fEJvW91OKF8yD8rGsGjmuI4m1M
WwLe5lztp1TdGiPOg+jpDrMsekVkAqmijCz/ZvTm0BML0f1Lhk6VauZJM3wfOClEmJMtHI+2aC18
EiNOvFFvf1d3sz4kqbKlHtEuVSM14VEc36SPq00859WQUNu3VsDyocXv3RBCikvsyyFvs4d178TF
3BjN9HM9LNjXkjCu/FWvJQFBJqfIVxcg280K4KRF1LBruv8DrVohmcmNFzIRn7qVPgwDG0k5x91S
TEQxoSaDnL/nuF5J3GNM4pyRKXoEeg2Q/4M5OdX0B8RgIJY04ELs99bEAaOY4W+xz9KTfaEF1cLB
tVS2WP2ZFYV3HJ1xd7VJXSY1+2uoJ77wnoBhR9jRplnwKP7bszr0yF6YWD7ub/NMzMByopGMwulV
ZAZ1dxCVZMvoe22Hn8OSQmEJ/8VYK0r3KsDI57vrDqwQfBK9Gc2d12yZZ/GFK5ug8YZiyCaleoGg
HpfFsGHT+0vPSsDXBAOV5awy1je9vYYSAxHygkxrF3H6apvjKqACGRisZSZQRx6BpGzxE83H4V9b
Ubc/tLzvTLxsADZXD95tpFN0GZ92Pg/nxsWr4CNyoKlQKIcixMZlvHnVDP2099DHqIjD5W7yiEAa
BowNw6SdxI24T/mOGvq6eaTl8ZzddfZyeyBhmpMnChOnqkBAPFgFBkqTMsSN8XiO0IAOxFCz1q3+
ngyLzy0kGbeOY0abiXiJijrXRLXBbP54Jex/qoJMIrORP/YC9pbM6ypZT8OkHidU5D/KxKbW2hIJ
50auU6XSoQ7OFO/gn4/GuMzZe/i/nNFMk+0NlYCZ6tpSCr9kls36rvt4aseQvBvmLf9IVw4IkH5A
ABvDxdfqDg4agsC4WMuJUz46S3bsnWkjISfXnQMXyH2tsoNREMtF/H/U5gjCAXk9Fwu/xjZ5B0zA
Zy6ROiL5WfxDX1VEyCu/yIZ1zqf3lV4m+3ru6k8Q/DiJt6C6HYPJLxKz2DcAuVV7SpineBX8hVV0
NsDDFDNp9b4Qq3c0IYfD4XsYuk88hmIa5POkadSEeQeRRNxWH7O6S7zTdJ9f8PDh0680K/wBVcP8
AoLuFI/DTa7GkpfGRubzlKg1nBa/bF+YB608aCrcgKtmcWgD+1enx0jnZ/YWowndDRrJN/sgWDyc
4haHBRBvDWx+tLRbPK7i05OkK7bEc55f60NMufFqN4NGD4xMTsbwxVL4qR8mA6rmu8VtYshaK+75
75KAMb7Zy0MyxZ7ma3JN65BJLxrG9R80Q9bRGY40qfQuyirQzik4V9oSuQIpSkRWb2dgTCk20OpR
kdo8/fRqQZds3THS6jqhp4GEir85WjyvAvVpCK5vKwYfLbiGLZTQXSV8N3Xwu7YMQHd+Vn0ciKv7
sZbckEqeqyo5rKgYqgr+n1A67bZWJgNQjIGEvx/CRKRrsghacFgEuRTm2d54tDjb7+6X8vlPuHBz
FTLeK5egc1dBdzXizncMb5QtL3NoG3JPgoFtZXQ+K4Fg9aFnKZqaKRXJI2yBuZzq6qdtphh1A4Ui
36VwYrOLivECIShO4cTw2xMBAXDE2XxxxMXcRjG79a8cc54yb1mbWmjIRA2HJfRIy0IJUSdCpOiN
WhKo9ZYp+r2Nsnoem8bGTIPcI7WB56PwIzf5unjst/6YBbT+v717t9B0Yh1gZmJNhpBr6MK6ixGo
GOjiNnmq2uLu24vNNn03lzKK5dw8AenbNV3SXioIuhqaTpNlPPtqNK1Q+xfgJibUH4oX/h3GCIV+
3WrGiwOBQcchaIt2imCvKaxAtxv3BLbFsh78cSW5xR3FOCGIyaB7XAHLbsgUczfIKnKJul04xbZq
emHW/DUdXBQvXnFuSSPluv1rVUUScr0yx812aG7+dzi8SxxraNtt5gGn0kePJ07OKA72+sts6+do
y/TWOvqqZy1JePCCXI5yJOREla1uP4LW/JUYDiQ/dYUh9Ze2MzEN+Cm7Mzh05xBFcQFcpzok8XdL
G0hauJUnsoOT0q++kQ1JKPw0dErVOS3JdnBYlVHr+TkB+Yg6GW7ShPYz5u+65X9TT4LxDekc7XCk
0AlA89ucchw362NzHCs5gu1eMziD+F0uE1ByPtX258m2ImsBCyPAE6dB8vDT9xbPDLGmTwIvPxYl
yTSEJwE+93SlXZuL/4ycB9eJ8aucMLp8gWEtLQytvm2HaHw47GzjnPh+miA2BIRKehblj6VHe/80
eA05VVDW/VzaW/1XZ8ayD6zbT8Lzg/SotvHEfa60HPoRcdwOg9gJHA0vOu8tjW9kgxn5J2VIoBJw
VajSk3biwL2JrrejdjXR1E/iEQImLFakmPlkSexq01Pc6NNRyWkPcPXLINYIjqdB5tORruN7pfD+
1kLDrs8tUvgg0leOolmpg/NcDnq1rDUVY5FwIZsLvrb0rcPiJeAwvIRoH/9D0txPcDjXMx47J2uV
2wX4GFzAhh3GKYBHR4hvu6Fhtu9lTp+NbALefnRCgYdzqpyvj8kRVnlzh8kp7rD8/bKv1eYnq9jZ
raXPEcFk2d7i2CNRY8azaAElEWlMUMoI47Me5bmdNakZTVakcK0mTLlc3+qTSH7FuCOAjxyZ+YOe
KQJaayKZIhKZlTOaYIf93egHW+wQKd16ye5qiIRg6u1n6jJ08VIp2Vj5PECHlwj6Wgwo4/eklc7o
Y1JFKHul3jtcCqim7ySZqf1iStArC+vQkRZ5OqyGjPZM2q/Hlt739Wj17KQO2S0fB4dJHdiDKJ2c
syWGNC6YhT9l+0wy9gCMtG57429x1DMFKEzblwYW45In04fHne/+R8uNibXCaf2HMzha039wNPBx
21conytUUYmrbO3Z6XDeCS+esZLMDYnayJrq/tRXaHi7ztapqxZ5gXHHwKXuYyINVHUrGGSVTBIV
87hbdf+m9b0MTgHvmyT8XtM316VqFpkPz7IdgPeLKRpbIQmORh24TGn8tDbWPFg0j9TJZFYtMdZt
m3NHeqJD8HXSdqIz7Pw1+dSW0BXU2JYpY+TEv/Of2hT2Sz+atlFOGGRflw9P7GVCG0nV4XpRSEuD
GAiumO3WD0x1hzPZL/tyUoFOBK1UPs8TuCqWt2TK/7vMEmADmANNDgRiWGY38pf3pqjrg8U/Wd03
EZxb6Q9bnyaOsUUWNB0DNOgPDAxozLH/VSjvsqVYE7ghhypS0AuceJWz8Z02cw2e8ysL+sFjU+Ye
ToRoMrKf0fzn14b3IZwHHd0se4Tz9nMnU0CL4dYtMsjhFrqJxDJv5QcNUf6RcTp4SL99Z8gmFjku
zjsBaWkJdIB9/pjXYgbW8mov3aNfc6ejkYLprOVBJZ+IcPk397itooH7X07YJBBMJcr8HDk11GYH
gld2w2hDtOV3XU0oavVYOfMliQUX4EJA/P9euetgcCKkDNkZ+nAdAUiburdH+VHV/UEVbYABYRaM
u+Ne7FLd7zhJnPRa7Ox0he5zoPmWnhPBtDyyELEVxVzyMSchD+FJTwM0EqjloSPwdtcAjRKSscYM
wgfd5bSOYQMueTpVPuRMUZ+2yf468j8kCcaT8GwAGCoyVtj81GUSFv6UCJ+BZKG4tkfAXlWGhT58
RYPdlBd/oyqbAFCc32QJIzlDGeLBxDf3mfAHV/Ihpq5AbIk2x3ObuhIni7XCsJpbEgGXBKmMizo3
JUc9168O6QHaAhxKMi1965fs51pxdukKz8KgtoDnvZ1X53BKisDmVGF1o24o7CHGbni4KIhgWsb7
1/7uHzvXRaK+EjIQwOpVFCvSllszb98jeyHBNpR3WX8D9zwmA+rv9A0DTUM0hBfvQnKmYVcWBWgx
HU7FvHuekVSLnKVPR9Y+xUZbI+dLmjvHyqicU2fZf1rT071SSyIy6idV7gSTwokSWi6PwO3Yd2Ug
GncrB3W8xa5QAx4Y9O8mrb7cjSc3mxgvdyNJ6o8zeMe3zFna43G+xheAm1iDpLEDqtu/jifKYGbp
cUM2EsWrjEyxsNcCTRp3mhKevWAlzf6/70zz62GVUAu/WeprWGmDyUkpiqb7QVK3xHzqU7qHV43C
6udimS5EIhqamMn1iu2JUKXd1UdQcAZgRQKV9jDawka7WDP5OP+av9k+hqs/9IJBMG/ITTNNsUaR
2++ewCndwpdeOBwaJ57JY16WQ5mtxTRl7Wdmd59tVH5ZznKUKQiX6Id1v7/Q9UoAH1FKSazKcyu5
VC8OzFeKTGbNbesOau8BM2PpE72b8TqHQ9/4y985aO7pIXCK9D4pRxSgiPtEFHsRP7KBaoLBBslL
1mr25rkAAW54fZNqcMoP8YL+4lWSIk3NbvMJSsnJAHIWfoZgbOwUeXoL/4qs4YbGJ1brK2X9s3aL
CFDwlMPOSUJWNLAtyLayf+jXLrm90fMjq/k2H9ZIR+t4LnFS+s927wJn4z8xEXIElQtjAGtoeu0e
4PJMIhoGAvtfmK2/SGDPHybP7pkO0CjB52QJCn7sGNvZ8oSkwd4vTJHbG7w/owjPJ1pfS3cuMlYe
/j1OA1dC3+A+7ApA16Aear9GxNCOJTM/PzGxttZkNnepI2wZnyMRHqTFcRfZ5+5tCozG/ucBsKiN
jHOxhQNPjvb+POETZtVYxpS5zXMldcC5BGb9+KEJzaQrn7tA0fWpi/HTRR7cjYCg0fnStTAWFsfL
MJvfa3+S/NzUpOlKVsa8A/aa+BFdYUSJjCZzEp9L5nZlJIAp0LZsBDTZMPxSbbIvePPLnqZqrHkA
pynkqUN5R2f/0UP9Wsf8VUp0Sl+e5tA+W8vSqWt7GSbr8eQI2JNNFxGO1fok+2Rq0Ag5RzY5wPAs
tKn2AdwyB+xR6+YthAADbsZNm2V+M3sYeAt/ZP4uzdbDqr6XowwrgMSJEFyE7L8XJ899NgcW9aS6
CZEPliiudsZ2jI0A5SkvLTF81mmvbL2DCLl8NS3YKewezu+haYVL7Qx0MceRlKoYnNewv8ZHGFup
EV8bS6hzmu8POdMVKHygo42JO5HW89uNjg4p06eH8HAiBB6U8z5zk5WKF0E7Li9ZG9Bc/HVISp+o
I+yX/bDmLm1kRzws64OdSbU+oJ6+OY7qaxrgJ8bOoncJOYkqyUQ2KyUDfltaRKQ93ahqF0TjlBvO
jlxbISrS9xSOiHmoIqS2Vm+UGWWiXyOhReY98V2u+1GtazZ3Rf1aAu7YwS/nFhwHXZY39g1nx2le
W94feCjphYsHNFaAQ/T6QO7t/0TnNH0dRo7yD+7wHEckT3JMlC5M8B6GpHTZD+cW7nfHdHnZqXYr
rZXZVr9FHadYczBu+rdStUVrg96EIW1ssGYlk4gVle2LuySceH6nB5gq1FBL9/qGqpdawBFYaZuC
GQaw7bweuvgqk47yo+0FN2OhoIwTlTFfV2pH21pX/qZeD9IuI4yeF1xab1NpXRIPH6m9kKdS482k
Y+OCDkY+HSeUkMeAt63UkgKi3APVHeDGrW7IegbJEcyqVe2TQFG+SVeT4oDk0WlP4nNXkHnavF/N
dIdSbhXKM47gRKPmeeXbHeAiT7jauBknHWdYxnjbiFwSNklt/gArwG/XifdDXEzxB041Emy9Gafv
Tqfh9e47dlr6A09hbIDvJoGVqfEsxr2QGM1Fsa1m8OtD9UGB9u1V3jpzwdQMzXC1lXRQQkxyk51t
1UMDA9TfRV8gyb5m4hp2O3zuwFIflIfh5AaJASH9t6cHUTkzwTC7xQ60iqroftpgmBE4x2VDRtUZ
ruVAfZym6C2CmdcfZrog0EeeQXxSE1z4lntFBIOHE6WZAx8/I1k2GAC10Cj9ZmZS6igMjZcPyvAQ
/0WptAP8IjP9qf45ALToAD/EThJvM3WDc5KpEc4v+0sFxnEL2r61HOYj1IqhtfmmUWGAqFJyWfK7
bjTZpzjCKDPOFnSPIciAlxx4wmUP7xi8vjiR3ePTcoM+BDMNC8mtYaw+vDmugMOLnPYzWE6oqrhS
hSlU2oy+vvu8uNDOQ5bO07Dp3XiESLnOnbV0xi48x1+8QcwOyV69uH4k1ouZUvSR/6V5vUG97CWH
EoYKlwOe/T+X6UzeAKiM0ufmEcJVK2bZX5JdLSw/+PVhVWh4QPIh+n1tWtvHah4dmZlRjI9pJt4N
N2U/SMisiA5BMXFX8A1hmLrUo77F3cKJhVp0V7tr38eyTCvcpxSEDgYeoXlnj8piXiEtodcRwxr8
pLDe/MJsA8IO+kUrnZdyeWUMXve/Oj5/MA2FY3bo7NaWNN6Enf/CsfyUarzxIlqxfvO4gHA9XE9d
Azw71DbN1ZeUithaaYfndj3JxF5kwU+A7u3h8bQgHfxy5eMZ0Umc6Vgsdy9O4QcJPUrFU4Y7HhBl
MrIRm98DuasZR81PtXOrm0wrDfol9HXTuZtHCoCrmzckyE7sKPZPcDertuBm1+mlFN2UsOUh0Opt
DFqvLrc3jOyd86jCwb+4AbDziHdkjB/Z6Ooi0hQti9wkYh0Ug0epuep/9nfvmXB+KBDaiLXzOiQk
X4UCp19lJXyyg/qYEZKNuh0WJMUtU5W+LgoWNqmXYZRK0OYN4IGL25M4FBSbCk5yKxRCcqk5RHew
xaye82l1gM8eMZWQUQlRLoqFuhUVgivCpGYJ94aIZRehc6/Lm+LeLT8NVDW99i+vTDgWQXuLYsMU
jX6lb+e8HuhmHWOZTMq6sflTBANFXxuvNL/uCpDAUXBJBGybDY3wwcMXrB/YMESGLIc7wU47KvVf
q5jF4ZvEs4PSmP6tWnuAQDc36LAiVMPZfkanBKoZdtCsxKBHx3ibrhi6Nl4SFh4C7+w+dA8yp9GM
RTQafFQVbbIFxmfZ+NKXIIS+O9JFocKzjdseTEYvno3loKiC2f3ZmxE57LLFUkYoqsCXW7IFMd3r
d0k0hj3MY+AmcJtDP8sFg1r2HslRHsj7ElV0b/YMO4XaYpKzt1OkJcFY1bThO/6XOmBuGMB4nmbv
Zx5MAZ+yMM35hT3bZlKymVIW1a9RTWhqmlNEDAfDKLxdqcfZ9CrUOpC7RM6PJdxBzRQmaB445GwR
Ct8vFI++Z4UlljKoR6qe9HxgPLjqDU4FGM+pEEwsgYFty6pLjh/1vGfb6mtA9gpsuXclKwAJgQRP
TbNYeLSAVsbvFmSog04H0CXHwDBxrJp8q9qdH+wyHjivfbotk31cibHv9CamiSujTnTJ4mB0WDK3
G76xW7CAj+Z5nqFPWxtXJ8I94rc9Ck29UdUkLY+cJqJ9tGvUoCN3bll0E8iHzGxBvqlQVcU89mu6
de2VuO5bSOG0cHGxX6QAHId7FPfYHmUPQUmG9nudlGO/jrtJKnoz14+ZWi3bLJJRIixwRUZUol2Y
HXJFL4+GI1d7TLf5SkHMzCYMwrUhj+AfKGGgX4S6sUiFwzdxAQZnhiVu9IuDaIi6XjwL6KrbImG0
Wyoo9ESV1JVYzxln1j/wQIB0oyHRIpCIRorETwZUB3FJxaA17QIH6A8CBGJYWFSl4XqxxcNOglFN
hulNOPQx/wS7/a1Rj3XH3uEAQfaEf7v/zqlMBldRIl4n1JAj0IT0gzkGtPz9fFoXciFQB0yyyxVM
JtVpgcEiHWl/qycclRUhdQzMwTI2vjNj6ZnqrpgY/taUVpt+Sbf/q98fOBDWivYLZjWQPZ6vOuzk
OtkiFvkI92xGGMihHeyJ+3Gs1lZ1csfktPU+spnYhxp7eCHIWlKyHgojTqgO3CW/QoSIkt3+0loX
h/SbjJCsBSamgBs7LE67LPrjzNa9DjGd0+YyMqXnz4dNWqGHJ7yZFUuxeuCiKYq9AtyxaJBFKPZD
nv4Kz5TTU0VC2N1vkklLICnblGYsKDrM5rfqgBxG5wnCHICFoRnGxZziYnkUv+47/cYM1txYbHSu
qlfqW1vag2w3D+9ve8Mkl2p4iXET1/61kPXKyBRBJC9lzHpFTo5L8DLwp8jrRbQEG6WU3lpkpQXv
5434kWQOkNUOx2WWBntLkxsAYMReNrKgCzd8INgcE4gW+qlmJD4EiyTW19c5M/bX+2eLTimA3WVw
c+Pt2PEl0xVmZajgHyjzddkx6ZANprYYnCbIfj7d5/IU272IX6IAywYNB2ycqLHYvaPFluNY2tuD
7ZwDuonj5qWuF0lD86iLsJ4p2GMVIqZQnKY0j3czck+YezCOKNTcki+TGqqRkOJ0B7vfzZTse4vp
bOMrfm/sl0KcqpJOYqBl+NLZwS37Fk+9muB7zM+5beCLxNWUTOkNbE/0YjYsSN2Mr1tiCJz14+KB
faC1jFW68uHrHaOQIZHL/b7qsi3zVd8UIz/0l5K+pkbNVK/0Eate1UAo88V2picxsKv9bG6JjUNx
uaa7EZe1bRyYePBohqYnabpe7PIxudp5RCRjtTrqxG5OgsStWXlVcayPKozy4HN36TbzY4sYg+XI
LGYnJ8ALgGrOVXDD1sj/BJYgBxp5BwQk078/rfpNywcLR0QsqdK8xfoXIqR0lqcN+mE4YsnbZwMf
tfHeMcQUxUtDaeS88dYie4qcnTvgZQrD92z6FuG+u+ydtRgtE0eiLbKUTg5FLpXQBPbl26Fgheig
CXd9kkZo+7zLp9NRiNyEJv9lTJ9YZtqSpnoasVt2GRGD5+cN2YtPXiyUyYeIt36Fa6GqCZgBj6sn
gp7zs2GhooKIW+QRm3uo/X+uBcbhKynHYF1tQZTxeZo7gKJETsFhuyub9HUoSWLigcD5K6/25STJ
b4JvyNXqJRILixyCfw92IkOMawgaq1KmEiyCdnj8zkrYwvV1X5BDaL5+ZKjWqZqnZR0NUKC6N2hr
16jiHMvyqZAG1Dnlo8/Nw8EL5FRtqtaZeGKtQ/URCe5jXXLxgfxDN5DPrAuogIb0rSzkOL+LWWmr
uPBZNpnjvNl5x5vCe37TWXkox1vJV7GGRRdRUVpJ87b3YBEFF27Wa/GMtgjCBTooKc6BXkyKI6zd
iO/dBWC9wsaABO+1nK6QIuRTuINm4T5En0tXwMgAk/AimjUXnJUNGps+HcHt4tIZhHf8hYFviA94
q00mvOuzuqnf+g1hPreZ0YrVWa9Yiwmxb7V5aDnkOjg2hf95Wbp4OdqrB758+cTJPl8LJDnd+fsz
KALweTCJpC1uKKFR+t510w3kTL5DOINIvdaSV57n2faLKItcfPrcmp3/dt/j4BuPJzr+DsqE6Wy/
pDgbD1jT/lFd2BhhgCi/wPZTmpv/Sa96EdwL/gSxjhj+QR6FcG7ppeOpT/vr/ajNkypaP9V2pgvk
qcmHDAWVmE9cJnC60Iph6BRvAHGBXP2+kVcy+Fh+mxWOa6gMC+gmIKLisAKnSur8H7JmbL6VBxaQ
/BvzVaHe2Dl6h4BJ7ALLNTQylfYGB1bPE25qOQnqZSqcibtnOSzUbhOoaXfWyPKm+aQAVwB6cCIq
jfU6fBfaRi7/ZN4GkWufH1o3vKeeHNclUanE315fSe/QwuN0EG3LsFRN0CdK3MA8l4zjB0n08car
3Kwcm4mNwbPQCX1ybNLYJi2bCmic7+E96IokKx/NiQj9B52mcFBERbzragLv14HxwXq0XfVm8EKx
xjpCxqpzvKoQFJINV+lLQ/f+MxuFptdqjtjD+z76T+Zz7GFFjESklXA9neg9ZACtfeFBeDXR5xr7
K4YUUiwdDetEo7VvtgH5pucsRytnLkIJnDdQBBbCp4xnn7TD3NviG7PDy8qyuEb7lV2ppivoKuAd
Ohs90BmI8FJY7P7ozvqSBLVE1b+75IxCLrUiyX9r8xhE1cIG84wmc0eOeMs413Zbiocsa1OmHjAN
dObyPqlSM9tPVL+/a/IkTJ1u/6nFkS2BlWKBLsPkGCGBjU4v0ONKP/5aqmSxiG4CUw9x6x244ECs
vOqPwO78gci5b22xRwrcG4GlJp1mNAg9RhbJ7V5G1BggOu3qYgMvKi+CPPMHvEwsnfbgs1YcpuTa
TcinLmbPHV0yBWOzBoV+PR5kD3hJ/+dxyT8ZMxynXVvmEToUYe40KmQ1hKcrId/fTRD0khJxu9XZ
OwiKq2+TPgXA3N53PSrv3JQrqf4IeEHRaTy4GypDkuJZjtFXTDU1DD2CybhiGoTH4Q9FV+Rcjqxo
gJSzOi0525SYDX8jn+V++Lyk75mbzfufgL6d09nICEvVIIcw1mnErR3VjjG0zw2AYkopwSRlToKg
Z+x/QTL9wrWPp7/SzLiAHLTZksGOXEHT8Y1k8ntZE4Es26nVjSGDxytW1kqPQOTAbVYSKOmsTBna
v9TGYr161AF36RwSkA9Bsz9qmoSnwIYnhLqHppw/05o8s3MyCBBk8unvVYtl3jYf/54l39A6t4OL
6MyCoe7G/++mDqw7vhFUGMzDtBxpA207vLIhQlmoTqCkhyYMoZuyu0SeIRuRhTC/SJYdGth7Nwjj
cunAjDOA8LO2k/RfwD53P4/D79kC3Hn1jqt8Whtjtnq+5tnby3UxDbDyHMSLmtbIe8finHhk3yj8
icXTfkJdOju620hEQp+fvJiunDGDRAZKVrDcZx4jTGmLAV0lUOV0FkjHJ++TEkMBRcNUKXC+BMnq
v4sLf0uVq+Ck5sVD2OsINjJu7k+COQ+AgPpoHtUTu1NXDm5qrbUxbxhMFNSGgbnqA55gFz4RHCIc
xqwxhl/Gy6qryGS4chNlF04zPvwtFv90BZDNkbbDbdRL8MKGeulVgv7FAPLG4TqQKjgsU4c2G7JS
oiUYWkpa3p0U2q/cKyujy55+y4BS2uXC2xpj1u9oFasYex3J4CGOdWcmIUL6m/nVi6c3mUE5vTvF
zTLfogiWFpG/Dq5ekct1fMjwuHFODA/qNXW6UA5yj8qLpcL/r3qlNdyZLmLRZEC5jo1Q150nv/3A
LiUCYIkDurqWS2dRh1umG8Bv6oBBlGm4DFYKrM1MgqJbqJkO/C6yjKrt2g77lxsSEHUDAqU29znd
GyXmsjSvG7RGhCc3/ecxt3k9gYO1aA/TcxtMriSWukseJLc38n9YbAAMQzbNpefrF4ELpsmp6AiI
6Mm2qW+VQGWp+opIjYsEtVxJ3aZ+Y4w/dpfUVTgJr1/Srm14JaoWHtbsLnRXn81fj/x6vFdJ+ZfX
TD0xd+PZy2aMu1VVD3PkRvJ7Jk67BmUvLWJLY4y+xKvnCS2Q7Ilc3rDix13TSFOeozko3aQrCWc6
suAa7COUzEMwBbjq0XLOJT6nYUD0JpQnUgneklUQGaydTS4A+pilkURdp1R+Jsh2GACLjBx9UrZC
Zpf1uwzaZCoOCslBPMeMWpEC4SJ0CgManLu0tV/j9ugJ06Nh7JFGld3LTwJ/tPIvANJ5v93pLWHE
J+xndEij21GIsR/Whh3C0samVnL7UgJHhVfnxA//7My6gmwXzaPJ8AVl25oaqK3rob3x0SlaHoRj
D+1TlSOddnQm56Y7dVMtXL06TkTQibfcN9HcQvi/PmuAYd67h6uaETf5FDi1h6CeTOf2NvUXltJb
jbQB5ZeDBq3x8p2eop+sgQnXJ+FyL6wf/wkdOamNB53jknNBv7MOed3BTavZEbuRX6BuqvUUxDLs
ZgUPqcehRn8PuAIdx3H8dkVx8x5ZPf9g72hIEG17N3Js6WbKoZr0zC273SatdEab+2UKOs+iNhfC
Qop4jQtyIG6nyOI4dZREcyfEm6Z0pP3RdXHFO/287xiM2QbD98qX/mUDYW9WYDFifQNS64yARuzt
hLXMyToxAUwjf+Z5O0mqNizTFS6K3QN/quY+4xhxH6tKKg6dJX8bzahPrkruN2DRv0f8aODA2iRU
sbIVjhIUfGpan/3cHHgSJp1xEcEgddO0WyGyN5HM06RGa/iR5ZvKC4j/UvpOkR6u0hbYftDe1YsE
ce3fEOwErGqgkSZIOA4g2dfXDnUhLkNrE9S67Tc+hmJ1BVhfYMyPaAkn4LPdlDTMbXrJJ4z53Y3H
XN33QQXe9B/CSUYwi4vGCSh8XyILMMEKsGXqYGL6gVjeLSzUGTerZtnsAEiHJdVVezQZN4CB7vPY
5/Pn6q7HhH+qJsXiZDE9detE6KwYr3YwYGas7UaSfDenQL8N00XS3qAysBjbT+DvJWwVxkjkYPWf
zsldi1M5hxpvfBUDcelyjhcouI5koTM59pe+kJP4bxdttj3n+XBpif9g6ATbfi3XhMcR4Uv+Wgku
iPUBBiMaofKT4HoITpC+s+0S4guPqLMgHooRrVEVKklbYmBKfeZL38ZApmRF5YTUIvnmhuomcGQp
pyGjFQ8xUg/rINPbmqVfSFiNgdgxSpkE6TXSaLgs7EcwnxkrSjL5tOCgoe/+TysVVYmAw1l4nTZk
ovrPhYcMOvpEVePuDnL11mDCdCrMYyCEv4c7X60LK8MQaWFUkEYPUXExAfz1Y+Dms1NecD0ICTw0
0b99JDa4Dw9F2OjCu/+isUFjXs9xmzvpdI4L0SvoLe5y7mBpM0vxJBExRayp2a5SGnAF9Jh4yFI3
ttqZijuHqM4YGnRAl67eGAKtfadBXcPpSJtzzFwQh12NDY94Feym9AO0WQrSsN7UMKQfp0d2nQ1z
JQqeuvm5i+GC9JRD6VkDVC8yU02vkuzfwuv5SKCTX02+K2gpNigzlokvSaLxBnzfP0/eF0cdttSM
Rm5rGuf/0F7NHqh0szQYKRqvtpG1zd0hNRbNiiEWogCHHv0WZJaQO3sfdOL6lwUHzxFCvn0241Rz
MefFcKwhEN5FhPc1Uvlhyos8T1b2WgX22LPqIujEqiwyKBiRvSsoRr/fyRe8/g0EPT80NtcmuAOd
IoGpNeBw1pq1EzLLgMafV17z1QR+/PPI5YPeMH/UwQXIaUnw6Ru7KdW9XrF1aCsUB5K/jVgdtb+u
xGM//sPB4xKclE4DbdQuo2i/FyY2kADuRgctgu2gdX8ASS1UT45kdPEAqnb6gPSnHodlkBVOI8pq
ZpHUVqWWIIUMYld42dhBzwd1Hl4YskEwHXDfu0HkOiN6yt2kKChF9gxw33U89FJtpQJcslPndMHK
ei7XEqlbl1F+lQx/gDzU6jUvv571PJDc7sTfZI/HQ2bK5i9vG75QQzuN4q1SH5KdpnT+RyKD2ydK
JskT3JHfkinvaMp6heucjat1lk5tZvGts+9pqroxfMOdhqUd6TPElRBTXDsh6OGlUDs2IRUH9uoI
uKKz1KWNVkJEnGTajzxddDyBiiGAeFnzRCOv5bgkoQsdJz7Fz6tPXFmX4AnCCJhnwDNQtPnwaHVq
paANspyQ6sGnliESC+eNJ9K944oM76i9NzjYB8D34aAUYazXb2asu0H2wVkSHSxiLn9UF8VVHbFN
cU+MIuvUUq9xzKqfac4QukwlGqjl6tR4Ik01W/z8cI1V1c69vI/BaWecOer2BdpIs+H85gfv4bjB
+9oKnod+z7DMVzuCp2aUcp3KYXEkx70xLa6vBQgmIXBEfNg9Ga+O9iOpy6S1LjOQMUxez1rQvBuv
SQwDxe/MHQNsIqVSAJ1sfWqRhKTfipUN576yUjc6RFNV9m+FB65ZUUkzEjuPSJdryRJ3dt0jTtnc
ESmPayQ/0Z1KqmoVg8UIAnqc0WCL5GS7jWcpjNlt7RZpWRxjbCFsoTBQro56ee3OSCO8eMqI2t2i
29RiS/P+e9JE119v0UvXpV4KpNlDTQqVIMqwqVaFiit56c/Ivfc+sfLaQ9tGGf+CHMKXEUxeCUEc
7fh/LEiDIscFK6SXDtPT4iWgyQJCXyWrfsLO1KLMppYA6EYXJpUDLnOx6sZzf0OF654bC1GNZhBj
Uel4i5xa8RT0I6yMsu2Ff6x5tnQGZgeM5TXGbsm6RNMMVhCNs+XDFv0DK985En1S+rMs2DDojLYf
0gMYQGQgREUYEB6ua1ZvwxsUNo2queVWyabmrEPTbix3SUGBhpxfPLHhxpQgUE7EeozWAN9T/2H2
hq+N4LqvntfA+RU3OMh5J+30WE2Ln6wvwRF+ZycSgQBpUAA9XTvcPBcAz0oLWHIvYoE1mFD/ybR3
RbUAlhfUnXy6B5skt005RCqDoLI2J1pazASFkDlbpSA9nP4J1hFa4/mmPTaY5V+y52D6rTmzCE40
I6ilZGQUpMqqt5MrTuBDhRmW9AI/h9JJZjYIpmrXpp9P8GG5N8osGPieXyxt3Dk9dOJcLFLT7eN+
FMALZd2ME34rKGxmQXBRkpWi+JLBKOnZ1f9QVO4dIHJ8WhTCS7QoD8V9HB7Xoceb6126MfPJNa94
2XyvdRDDlQwtG4rQBogMIGUJn2vDiMwIMSFolDYsbiJo2DMk9v7YVJGhzYmgb/UXOMl/0Z30lYSF
UgFiXQhVm3J0ukUWZGTdC3UAb5XTduJY1ARPKUa9mhaabXQuaVcHSUwOnfJw2uy74/YOOHu4f+wo
lRNFYuIKlgip7WkFMeY4hdzUPDljtyFXvBXz+cDysjx7jii31AaK1p3eVameiyv5rhO/4OSaEFHB
qcLfbct8zipH97gjPW30WD+N3l/AoDNa81Lz1bHvoo+jaqN4CoRFFTVfg7xgvST/VEHAtPbvx8Th
npuDzl9sCTqvWNCHabP/TQItPwIljVpXEy2fWQkunKiTyDlt/m2G9x1ikvpsc2qlo6uMOhkuZ7f9
BzZvcJ/zsZODyXlXKT2cEe5WuCFU8doqKJi58FhYD7INhwPS6hDwDF9Y/1K33FniV9JhXY823BDg
8UiNt8D79577uSpV5pL9lTRGbcFR0PCvX3f9VCj76JYCno6mS3B+leMUjMivJubCLWCQWD2BfsJF
5P0Wo81051F8SA8z/9O2w8V2YgbPXzuWPAjAzjhAUuF6vxcwRv94GjMMIAsDGSabpSJCZUavFHzf
q7AbNqEEGsHd+H7lvH8AMaWfXBjGGu3uRAZAFArfmlCyz5/3Ywv84UgzXKDFgrSlv4HLsQ7MdpN5
lJMn2oEF0FbaftorYt6F8B7alEr+QCykA0CrB1jZQ+30MzApQ2WY1ln47FXSyz+DpHxlD1nNYTvZ
JxY0svLT3jOANt5ZBYvC7UZTOUMQ161cGf/qH4ZKfHw8R3mCbSmUPSN8wdff88oyBKFx9e74kcKu
2S5x+dTfwnjkPGCXsFMaMInfxrYqpxaHQ65R0+mKPerhN8r8aill2BHZu3nzJYLCEShmOM4x1Rt8
PwbttqsgQsitEhG1ssejaUiafe2DLnei4OdnSbHrb2yFEakq3QYMd0WYoeHlSyKNNPGcZ26eT8B/
0gRu4r3eCFNYFWa6+nY4on+gFjOuQoAF5PyvrvssDq/gFUaRfRlZL1bK6T/g4+6nGvByR6gqNzKx
4gyvDxsyoiePrBSASmxnK87WLPrSGPleDZmIsKSK53qcLtl6bfcRR3+z/3jOfHboxv7zhi1KGWum
PiROzyvcO+5VkOEMlPVFmT6JPR6YD/+eLM2s6w5msFhde8dPHhDkwk1NWSkA/ACef7g5TIwwhKho
fRH6tzv2YJzZAlz9JjQ1JuV5FNL3hMaLEXlTLDtfOTvACXGBNpefOZlGAs8TJx/d50OIcQU+E1qM
7Bmb6/riD5DQTxfW47SfpwmwKj7jHyOiejnUmpmsx6Y7J6+PmVFfaAe9BdyaUeb5nwLWO8Qa+Um5
Ejj8vx8ia2yIt2MV3P6KfDHSdBw2xcUaSGXd0vF26SMEBjFacVdZFiiIVXyZNStmy/SaNW/FEOXt
qWaGNXEziAbwvD6zjsmWB+k5oXX7V+FFy2mHZ0UJaSSDv8V/9u15pnhojWTEoeGfk3nP61JIIbCY
UKEiZ6pSC/lskeghtSVdEe8LM/8Z0tmSdiV4WcXGyZwUDIzut2nAJnsNtqhG/zplLbQjAQz5YuA1
8GawdPLJ1WXF0uRql80Q5lFII5yOjeTrhDDdzaJjVzoc62cBOi3EGxBVspE38pyhabT04pf0noa/
39bdD0Ilk+jwmMRulOSzbPv88TMpi4my9UWCmk0fjqHhTmpAEkx5jZ96EoRkSt7jvJUdOlQb1toZ
n3iFJsszUVk7WW4mCOkEwJ+TbyM47kPaUyj7izbjqHAI7OFUU5ZJ7ZliT33rmN8klGakQ8BHpYmU
ruuZqLeL2kA5kwA6qpe7/7Y+nu7ciKWFVmYgib/YA9vtc3Rq5Y23Ivb6xyhp/RFK/H4d6pwiB+At
0eha7dZ7t2E47LTJpb1L125VjNKItneF6t7p3JL/DXkYDDsuhbjMjRLFrvu8ukallyNU/U7cEAk6
Z1c5fmzWGeCUn/ncvC1X+IatIdqtjIcn+Q36vmcx0bO4hczwNsSDKHmiOqCM7x+H3qiELSftg52N
6tizWzFqXLG3eZtQjx4vT+p1qYaXj1kqTUEN4QXX8A1Mh8f7fx+pwGSDqzjw/VXy/DGr2ZVb4ugD
DVPuMSNo46flEasmEJlb/0+G8dcukQOG4xTX8b/XTb/B2VC/UkBjxTfnmsyWP7y3QF1y7/Jn+37e
OT3JnSeueSKr4YL8QN9Im3c1ms2krQoi6KOw4zVpyGHmcGOPZUvYp89qBRCqQorx4JuFYxFldKYG
5IBh1yOFFZ0BZp6x0XosrGfHUkoravWl+Jzu0xzEjH9w7iKca1RblEf8dQsXP58JK6LNKyrYoTvp
BFec8mjeQH+d+NTqL/s47Fl+fSAkLK9zlGOsHvq6prrV0vIYMMUZhvoNz+7Tb24TITE8AhyyWj0G
10HCefeH3h+FXAB71hZTa21DQWJnWYlWfPbq2XbpsxRezXrkKb+OIPhkqOoB7gt0idZQkrLNioId
CQ0U4i1/7IUw/0Ueo7mGU3EJp9oYBuAm7iKaA9JzOiv7ArMTZm2gBaDtdzwTWmYZWq0NUNqyFoqO
GyFBkCqsKMCdnoGoT6UKt7IShHh5Uc2f9MuHN4DUt6GdjNN4qQTZo70UrChV9Zh8MqebdpWfPMq4
FPRIB0Lz6bRp8jj8Y1cRd3gMlrZHHaqjhL519lBm1OwvqGrEUZDySOI7bFHGvSwnXHR2AH+N12Zt
OCL5sto87Tc83e8vII+sGa6maDfzyYIdOCWcpgNOtwkQyZAJU5oVqQycDST7sQHCv4r06KMaWfyS
JqysWV+MIGZDG9rPTGRM2tljzDiySj4aR/ynIlgWAd/sf0vi3ose2hz9RFzHfxvZQQ9wRfGbBDy4
1GfPvTiHDcXXfxFM1oBXdRFPzvT/5FWGGQZFGf7iPDUW8tKcj+J0Zn+jOSWjjZVwieY4/xYgEXKG
EP+stYwamEZRajHeKkeW9t3fiMOTqEyBOmW8fN9hFOuDiAeMICXkne21GDiEYvHPbHK7ng5BmQC4
vQEg8O8LSmRAsFbURnjyIqBWe/xuG67EzHYWk9AqWt86vbu6feOxtwyoPx2fKMwXVdStnrlzxrdk
CKmJW6XCjpnbtR2ibjOwClWGW4c5L4FWPHS+mo8UyM6C7RB7VZ5rX7au5nyWjzfmvsDiu9cM66M2
r/X/i7TtGVS4S22g3/DphAutjLb4kcYxTLd9gcC3WeQAuC2ag8NKljVb8LvCCDKCdHV5ieXpYtkr
YgpVUmeBdAzuZM/ttmkJg/KaoTAD2USn/Z+HLal+9aMqVRQVdeeOkVmzu21e60NrMFqDws8tHxf5
9HsfracSBQKWrAHDLKekhrDc7HfFzkm3h0tyB+iKoUzHDDwk7eyqDxGz0wb3VzXpUs/TvTbeQ7Vk
BByvJQNr4i7+XGwICT26IS0IzYVer2dxl+7S5wEYXGaVIfR2buuo0IvZnUptB3QYYP2bCoggjM13
0uTr2BDhb9rSgyxvoDdRjccwjy8M8f0HbdIpxd5jcVLKn3bNBl0QVA+Q+K72rSMpinIBRVnSzvlJ
+TGLKOpxzZLRGV1xJuC3KMOMXAedIfsvB91B+l6UbooLcHgENKIY2/cK2GFsHyoLfzrFecUoV2ub
tJRK2mtC2Mb5LYxOOaKdoH5wu8Jv66096IEPOTOFDM/m8/efx382Rgp25Rg6ucLkZPlpRnXDHj9I
fEbjDd9OnSQqCVK0IN5dLNch7ximOB56dxJLEDsuN5AWn9wJPN43WBj0H/JLIUZcbklGm3JCQQP0
FxmbvrjnUr4xrkfEPfUeUYcDcAk1BDFhXTWJN1il5RtqY4WpymBZe/kxsc+JGPe4yyoSgUFJ3N4m
t2lIYABUVxeJzHtFMqrZIWFbYPKSomcPF7xJ21tu2Je76P7HnlB2wwMVr+4DGRZUHk3dIhSvu8iF
jtWLLEqloUcAe1Z6ftM5s82M00bSYowIuneXRo868GdkDVm17qIbaUVEND3+OrC43IGNNGhTcGH5
3T3WwMDTKblCo7brOINEcj/kDa+xx43Sgd/VPJoiK3/fj+dNTGULRI4TwwO5QNY6U6qhdLay2fSG
Dzh/kpSMVIcxu2bLcw4VTpn99ZcuCZmz0RWnwRUzKiFbXkJe26APjepaTvicrqOj10URj8tqPkt6
RvgEqoyf9JlelPbjH4W4rV+C5uVs2IVL1BIhxBrS354l4ImnOMWHkF/07mhtcjhe6mLfO4SE4YQO
naPmLPAvvE3sod3HAKMmT8h3r/F+IADmPw1Ab5HX9KOYDu78LSNgQGGPsVL7ejuP4jY9ExQnY3lU
SDA5czoqIiTPbYeaQBhLV0ZPUjphFpIWCf3g5FqOsDG3aKi/XFBs8lYhy0Zr2iKhpFLQDLhezg+H
hU4NauiVZSSf7KRmSatbTtru8DVq7AV1+vykn8Fe/afyIM0e4HhJ3E8PRGv6VVod34GX0Rdip9D8
MOP5L5n5lVOXWTBeterCn97FWUcfHZpKs2iQ95NffBCb4Ahf6RdzX8kUEOlb2s0/4fueQmtFSRON
AinQOp+bKImPxPim/XDXo3BsFkWV0xOMRpAD3QNRJkll5f/iMftYXYyUnf1zA1KOA7y3jSHZZHds
9JHCmU3YtctpEY8Aeok0aAcwoj5tmt/MKEQswnX4LJnWWcl3yy/7K6vNJ4pWk0JSP1BSQtvMkssq
6KQB0JSTnhcn2kxrMmMypqkTXJC5LLTt8ePq8z5GMSI8Fqek92NO26rVPRQ7Vm4WiGDho3YZOp1x
t3wCh4pUwh892U5Z4Ki5Pj5v8knqxZy0q9qcPpHMO1DjgqkZ/n77Xp6xo/TJQOaSg7npF/DCVF4y
34+zVOp/keiZDs3iDCFWqfRSpQQHmO3ck1UHCujNeqV7rdPqHSqWHQBRe2r1NFBm5+M4aypSsWWt
RWnu+tZdNTfgq1Adk6ZbEH/HmGYEJ+0Irm4bVunzn9kci8xw+AmTZaPTVKReOZtti9VVeDjXQjFC
Z58mr4NFIb9p40Wv7m0DKz+OcpLKMK+KhiPWTLBjcCUhWq5ZkWA5x01y+RsQ/4ZlD7y4VkdHgKss
pXRs8zw0K0i071iNawZRN4oV2+U7ZL6t1xEUfFIXRyphR/qXQpU8ojz7546LYCpFDvn2NEXk5CR4
Q2pPNQokXRrXwrXkDA4irOgSMHNXn/XqefG/VL1ZyHTIX+mirdM+dzLQTfmn0xk4UZVTpMlpI8S1
TrjDu3mTFx5fILLWMLYIVjz9X4y2QSD/jxup0IxWCRR6kF/KTxv2a+E3bX/1HBw39jSTx8xz6FzK
396r5TdCl1GMJzVQt8f13nU3r9xmmpmAn5Pt53Peyw+UyN6nvtkS+hbgpiFkfJYm/0BztXBDucnl
U3aXFVnLFVIbSBMMfTSUwy6fCkBH0WOXpGA+Azkgj3iYG3ZSTFhJGEy+KZjsWh7Q/U+nTbjfL60x
LtmcPLGGctbH5c848ae6BxzJ6fUmXuJnYRW9FZv9Dq7G91P/nor1ub9potTn71xPeROE+NvMcDD/
+otTTiqbsoIJ8sIrNKN8Hy9LO5imv8fuSD7dHRXQk0JDcRnI/GkRu0MwJ39YYwGY8/HXqSeMSgCt
Cv3V1yl0cCCpIwK49zqfuUTaIGEQPkeREA30IrKA8Gg8z5JcS69F0LP14WyDANtY89J+a5ZKj/VR
0vYXjOKHy4Gsu8g33svZGRHkiDVM0Zf80CBsCbq8ukc9mqPwsF7qfwlGHdrCHreq0m4/xWg86u3D
XgO73dhJ7ZmnlrKQv7RuWi7UsQ4B3lnk3hRZ4rDx1y+g468qCj5UY0HeMw54niV5hTYEvyIjbHfV
M4ATAgyORKBOOv/zkuxyqp3bZ4JyAPYNBe4yu37pwS9kTR5ZMSfNl6pQbOuqpcnuhlD2Tmaw/atU
e7LOZB8r73EPKv62yzWKMpd2enwhfdxmoP9Xh0ElSD2oGi9/9JlGh731+Hs5zPGijvHC0+/uMcCO
3yhc1NBrky2KjFSwcBCoKjxG1mzp/vY3b+YFvy5XTkRwfVyfaNJCCD0/geGs2tilhi49n8MWP6S8
lJLQvu1I22L9UzWT3L4W5WC2DwGh/zArssNRl4+wJ0VUq40/DVvbIUbjXl2b5j+hmr8p/CA80yL0
qbH6Un/1B287HYfbqFwBHGF9mlIkReyO/ZLZXFk4N3Htk9CmBZa7Ma6lpqBPkd5VY0T2plDYVu7c
gQZLg6RUG8XO6vIMVzNVVThwgdyzUqQ3rZ464rM6GUILyq0qODorRqSftZx9vIR6Y/fqkI314oBh
VpKWCP+m7WTxPrsCnAtqEKs0RWEmUmkqycUbH5BUtu3sczqH99ZpV3dWO+la4B8HRq2Q7GBT6AxU
DxB8soTfzZg+BevPenByVsVyKVn1W9Yf4V4VCYau/cLj0pE/m8pXKRZLK5ifhb6ng7V6Menx327s
7nL9LFjkpsLSebm80BTPjTI5vGSrJdE40SRxSrMgV7BzPpPj6Kws3z1fGOXKwYb4cr4P3REoDYi1
ToRvRHPpFaVrjSwfILKXrOPnAuJCL5pp1Dit5Uu/IfPi5QQY1FU8F4ymYajxw9AQW+U7wUGryg/q
NsBqzM8r6IONX44d5EjoiMCyUrJQJ0GcYL2JwS8UTn9RxidyiCNqJDPTiZihG3DzDFb73x8IUsh5
m4Tnf3W8EfGUJsF7XaIdOklZzgld6LGedQ/Z0emz1Kho0dsf3OrkrnokDN9Ey2AkC8gU2JBO7vMM
/f2CdWMKft/T8AQTxBc7Dp2VZTCTzGZfPXy2j35Ogm7upuWxzCgNGfW+eQwHTWZsZDVsG4y6r9Dx
k5pD0eF/b2DnFHE7wLMdtzdzcgAfm7cDUPyNcKP1dIbgpx4o8zZMXtcduWOdbrAX42VlT7TJzlL+
/0FRdGz7XZr6kgI/NH10bW6W+QSMK6PfjNMw2m/BVWO2gx1k+rD7A2qUJLGxBWwLC7FBP3NCnfe0
f9brOREpyR1cqa6U7Xt+LP8OxlArCluJfntNYE47LgWiORhtHfVYlzj4rztiQBZNSlrI+1d1Liex
d4hkJtRNFND13M31xlkZ90L3r1Gqnbg4UL9aMu3a54152+msEa6OXh6EGewTrKtKSbADaq4u0CIY
mbh6LROYD4uOb7ddjIdHtGuQYHgfIQkDr+8GlDz0sdsOUGTgK8fUx9XfhVgq9N+n0XfPjlTW1dsX
86LnFoop8CHvBVHGfmXqXWevfbOVBc3NN99M9tTBN/pSjaKEBzIBsazNOrjtAQf4vkXzF9MCmAbB
ORz+RXrT8I4XbP4OOWKuYjsieQZRJllrM3A/mgQi79cvULkOR9Ryc3J4L5BmdsvOURlc5r/8T15S
n3QdOuczWfcgxFgdP4V4KlwIpFePp3xF2aG6DS4YJE9te63Z59blAJZVi2peItlpFmQxNa0w85s0
vc2LQgnrwCW3ti0rMf3TABwoD6geq03D0U4t1YKlzNCdV8Cnh193iOGwMLHlfdVGiCjdTpKBMtfu
IWA6iwwqBNGgKRN/RT/CNRt+Vt1MJSekrp35Lt3LI/9KQzntDxdcCjv+oePTd8mB6XLnLLAchSTn
c6iWs9LqvMO2AzmUuTXZ1XBcfrXamb+TWACzs+6xapaHJI+e18Bd8EAP3FCINf4LerfzrrpRoG5B
36pPG8UQJza5j3dsHP3GgMIK/IcmP7YOh3/Rc+3lfgdaUfI/2tgqFCJVEAARijelCReEp2A0qaYP
WrSPH8QNJaRMLVK6Cuqs/mnEbr8uDI0bbW42U6dLEY3AlHKWq4c6oQnFbUan2RtBTKkbPVscfuWD
GLdcO7joy2tJbLiiQyzAxeQhaB6bFPJKfm7yfJxqTLB7x5M1LhebaxH+VvgLGRkGZHZxu0cCoC3U
jGl//RyNQt4fNPEnZ1V4cbRgWe6A53Vfo4AB/IBau01W1+YOzwxIvff4gMFUT8DJxZywzy4GwI9G
Ekflx8aXBj4q67Vrm7ITDAsQHl984WF41n6WYPWO86pCixkYm9c0WAVSaT/gfrgTxwOblCS43wyq
X0Qfxl322hpukIGo18Y46tX5CfUOjN2HVJHUCCGlPM6ssXp/nXR+qgl5ehEGzkcxLcVrmPjpk2X3
j+6OI4gPT6yIU4ZZ27fO5bbTVJYK7RzTQH/DAdmxKq9JFtZ18vIm6tKqsfLP/V4yTacjK3LG1uPS
45nc3M+vu5CNXlhvUNPylayks7WYBrMKld1rqW7fjyTwMZtG6gvwX2KN+Z9uE0g3kWX9vjuXdHH6
2yAhEsmrWqnXeWHk+zHT5ulPT9O1GwTWR34KhkqB5g+lGpMtfIeKXaHPizdGkVqccvn0+aeiRPTO
7TK/iepXWmU5INeWGZ7HOmjuBmAb3biOrFb4jk2fkPS0kFwT6A2v1M98DCfFYar/bMIrF4JCRZ8s
qSd7YwzVhoYI+mlLdC9jq0wKRM2ySTK5knEY7wBQNx/1W/wL+KY6xqsJjo/kAa5cWglDP4KM28Th
S8iqZiG6rac9mDB8KscYp+pKQsWQOAVvBUau54+BRKyFjD6M/LtL7wBLnpnjXYJUP8FNVJEE09yg
pgfHwdCWtJKbhVuncPnge9+ccIqy58izuacSnnyNETNWkQXRZRPqPEMy3CkpKpwrXVHKr0wJp544
+bggarprWysLdIv3CJ8cujKoHQGJlY6qyok47CoqhYQpf3OqnTSWVdzXgEl5CPkwM/cjzireXouJ
e/zcmJ91FXaLM1dOngd+flWGapWcwXCKmrPB5HVv9HEHJs+r8WVpRLhMmmBdLtIeEin4HVmUWAo/
dL7gsNCEF2WL/gND1lYNiVPkgNKPVzzpgxqKqu4iW7kacy56pm9ouMQyDLDlGiXcz8AvDFdBL40V
iY4oe3J/tVtdLBA2agVh0TPo1OPSyeW9G5xOiXYbm3QMhDl91eulG9psnkbWweqn1zx+eByNzUNR
NHSDDIgdHF7VYEfkdfuOSTOqMcLSZaXxLGXHYExoOFAgbmcSJUL713Hl6PYm3KKQN14IYvg1wvWQ
c3+l96nfiZ4/0xuxiERPYvytmbKIZIYBB+0pf7G3y4hmRF+zqBp56H2h/kDuKgDoZKPs4RpEoI9I
feiLkwMyOUNjzcww0BDslfBbfSVKXnR0N3NDprU9zOa9l2uhBk+khGqcemJn9Ik/LBt/2Yugq/S6
dzNlx3mSiPnyNIufS2LEtcEIrlrtK0CWcqJrjwXocClKruMmzCaZiUIjXAvTR0FwetS9TKyUztml
pWHhivK6NJfbKdMrGRtdw1zcO1wAgbDUH9qPq24c6i+gvhsGpOLrUUKVoX6K3umDRnS16OHibaYL
htiX00f+VQ8eS4xlrRxRWIZjX17rFcMYsoS0YZiLc+AFw4IVVDSrFIIme3c3pUlNgspcIwL2J5Or
TTh/9o5XP9I7zlMkP6iNHkLRXw/ULAawL+/FAdyd9pdfCwFCE/OBs0H8bGf6rjwpuUvx5D/yVZDI
FknxYnYWaAwR3Zdf6TYbg0c/jl5i4YkWoZHJGLSZWrvxQCkS72TJ3tmobnw5jqi2GAm37TzjfP1D
p/vBU/42WHXvOp85cQMGT/QK+uaalmpkXP7hQ4JWBhy8GQYONHGLzGPcPiU/HuFDXdtkIHJ8gshR
jAInTIHS5RDlQev/xodSV4CPtjfmZvL3NZ0RcQzyE65IpC3qqep03JI+gJV0EbwyNeSiu/lo+pta
5e9/0Bry1MDsxuUQdxD1jJcQXomSuJnW7tHSiTO6cDwBHwiqzFMSsSPWYAJ4Z3Kddj+ypPSNqQfQ
edxSV1i2qHesN6dWjjmszLwc5ZlP/gnPokfWJ8xl9vhK+6caleRk6VuBypTdJUSF3YtBvZIiQ5or
eft8dg2FfserRiYjRcS+d0azLaEJk5PHeutN263BHe0snAOIfL3RD+N9ca6xlfBTDjp69FZEmdJu
hcyxFJw0OVz6/pMWumm+wSEU2BUB7gBAYt99BtRnVKuyEN42D0dn+BkfM7Q2SqHQAbGoL3Ud34Va
6V0DSnmu/SQISyAIeiIn93qS5IAGv67/Df3Isrh/islgbO9zCP4MqFzGTeNmIlpF+ZA0v6naYPTQ
TT/KQgxPToKhVZ1cVPNd1RrMW45vLaxa9cibcktKBkGJm4IcSNtypDywth74XXk8FyzIvwf2JRZf
uqwtWYLH1W0rA/CPJnW1QC80WeuVd6zszg7DBLdDfssx2v6esZtwOlPOL8yw2h7ryB3Rb0efhV/g
J30YyPZSmZFMeMHgPZlndhgiXwC4+6gRGTvNmuy3V/UAsjo6y7NBQmWLac5m2AFkKIQ0X4S8rpz1
VNGgrH9O352shpeYjYHLXnzr0rwClfRHHTdhiObEczv6ndqMjQcA+OZNlwCrvxTnZOr5U+F02yV2
w/XkIsr8lacw9bMarfpsc1DWbpSQkT3rSDXtmWn4vATZXIauwdT7HzB5P8OH+lWOnhscBe4zCxfm
5iGNSC/wx/as9/RLUb8rvRUhlC8DUa8zoNqDjzoU6Nlt25IBLlDq6ZP/IwTuIC/w/OemLFUxG6at
PzOZXl/t+ODXUbFgO3WSfxzRuf0LMZxVWFMT1RjwZcNXmOoaRmkL98fdgsbZD5tUT2XRcx3K7XxQ
U4bPBgi6l7rr3d1QZNnQrVNu29n5eUEgTMTCDdad7QxYKr8T1Vruj3hnNWechKsYcypWxFCathqg
HwvPfW4ipobpn02m4IgpU174hrnmXLabE05gEJq5yWZztWJmR+TlpkbIe7yzuoIGJYSPpzrc3umH
1nDWJFjwIcXQvELABCsz473IZosdrEbp9TrylP5++wBnzAl+GqH8QaSizTbmBYVE9zacV0SzWamt
+o1zc9PVyKMA9uxzKo7I3xYt8dD1XftNf52pEXMxVXdYmYEj+eGIZCwFUWOa798QyIApNsFcFmji
WSIsHG9dJtcuye4u8/mtqzJMMSKxDOUfBIP/PGbmn9L96NBEv2hldJjEBPKs6IGTohq6A2ODenyi
+dPP5cFZ7X0r2GbiPCXT3INJmgvs+nbsJjeW/1rNBBZwMBA+nSxvg4THYW/Pcg7QGpqJsQDl8OVb
K4EvfnW1y/qiNMMZYJKw1mQKatre2MmRb8hQQ+ayaZqHKJM1Xbj5V6Jf2aO71EzihFLwM2YimiEa
JcZGilNxzBIr6NILg3/t8kQ3XGqie0hqlIb6JCVyeyraTerm1FfdxcL72yaZKtfX3skKaBJTx9M2
6wSJDWGFVwgUE+gkJmjt42oty1nonF8SsiIENL435cOcx3CBcQBUmiJchSnV07CtECUB/oRh+1gC
9+gu0xqiprgmL5ssftBnJqEA5T2iRsukBtVnXSendHvIbo1jqAcwTsVKCnqnTN9cgs42Y+jxK9D0
kNeWhj0dZczdLpfh5ZiOZlrfuigZ8bn+xilYsh+xSEcyKiIgegU1ThGkNbHpyEeUdIirCnobFro2
4O5tVvK/xPmY1XzKiGh2EKxU57ulxJqaovptDmSoRg9tuJWlZEZdBpImEjalbQ7FhiQMqEbyIXFY
J9zKTBmjLNJRxqwZQpkJG7Oi0AITiQlR/u+epLnxEqXv6l376H2aRNud3n+nM9/qMHdWAgMeua+E
sBnPxUwnwD7+uMWO5WWksFENWMjHdlKjeFlDie5l9YaccYZhc8TqdeuuVFvrZeizslDUA/6AusTr
KAU9ToRIRBjztKVp6+2f6+aM9kB/oLQW09772x+ILZZE89FDht/V4qVDnA2HnsaduXSwDU8TEIKm
vD+5IxslLUDqj1Xa5y9ZL0Ff2D6qgJ/5clEqWiSRy5mBDt4kTd8ZjFDoXO5PXB1loiLtr22RR4GV
pT6ZK1rDFZIBTPsUZuPGXjbNoTvSyaxd3kQ9iqiQiDHVHvj1Gu+6K5TLClySJpZ51JiJvnG7NS5c
dW3fm6p+Vb0b4DpjmW4/f1mODGNFeyzop7gB7/DqdF1RLVL642a5tXzTK4yib2CwwQa5agFWiH3C
0kLmbzIxRfKtucRg0bbcw7v8TTZuC52w1Yt9qrx2sChF4gvRT71ck5Nk1mdEp+FKAZvKN3w4wHZi
5aifWEU7R7WgGvSYu2HGWDUN23cUe2ltF7O8e85nTWIc67ZCqnWi/XazSXhFcv8IC+2yYRdEh27B
x7OM/CeuoIO8wwGtcL9sZQv3s61qk0sSnrow321Bzr5hQVHF8D3EHSBLxmuKQ2iZO9Vr9ffpwhiV
DG55uIoTrXJ3UGRd2eEH5x3oWscI9DIQwFZ9mWyMp+kqo7omLkgjqpj3A3o7snPnw4gQnW6L1Jtb
k2RLUaeVEmWVeQklpCO/QJuyb2/SGrtdADz2Yp4fX9HeZ6JFuyyE1/OhEFtlSJnND0TWvypzawGC
YN27xo3CfTa+iMinAxFzWuzZuQSqNDVdrF4boFHOQfKNMiIeJUCZ7J2a8xoC/cdYbmldlXeZeeYv
IFWpvWNOxUe9f19ONhl01pVAqk53pIzlZgBPOQNyFBCSTqRcYG+vu7IP5cGDJ6sBHu0ZEsosjZLX
M5zF3nAw2onH1BKrZrZy0Kt6p6kHsiS327vPCqNg1yV/1alJZvUoY+c6gr2itgM6uRNnJPMk2ZWc
bY634qvn8JOfWUEwhC61T4RUn2RLIhF8nTq4oGRd9LZ/5tPcIbyHzyBOYhUaW9axmQdu6j/2bGzH
ZvtMZBcMtYHQCkQg3e07YMIbxoeDtpUpNZ5xcyqzYEFPbEPzX+t+yRrQMfnBNUjJ6WnMaXV3ktil
5frosXOltWvfs8WANk/iIqdyC3NkHId3jO9gHTrmg+cThVvtGbjN7fyqGNDABhDmKacmZ16ABMtJ
V1ShFXhR2wgbczsB56jdmAYb4LVIAL/K6sIVtOAXyGBmgZHu4Hq30q3zNm908fXO5Gqcn+hieVGW
Mxp6tIkCoefMrUjaKt67AeK/kzJmCILaw4DZUu+8NLJovEmq6MHifst0iUtOvETJXZdZbNl0rsrL
fRtw9RRNtd21l0m3B7rc5x6a3loEKZQ2qw0hbtc1fvOykyYPTg0r6XgjV+LK2AUyMHRSyayCl3gn
GHMpwJPzszIfBswEpG28qoANi1ZujId8rZyUcosPjNd1TOsNpJcNR3qLrTV2Tp4K07d6sDlx/e7C
QhAVBL1TpoSRNI9Nvyzo3o86hVveL6uWqxeKjK2spJmo3c0jz4ZL5WySF+liGF0WZejLaiKBxdfe
bSxc2Q+Ur+kEbDNjBBb9QFhrZDkzTliUE6W41QQ3/ThbKeSxpcMP8PgSm4yStgLfkqC9hlbhqiGD
vk4lFagU3Pt3CN7nC3bfIzi7D30EbrMBBtqjdjFchEYPFdmExmgaXDwUs93xyQ+1w8Rr/SoDOQdo
Hd0YG3J2/CKm/rOf14/9SC1c+VsXy/zMkj5TdxsTjnTIbNjqAwIyxwSQ3V0w4N+s7Iq694hqq2H1
Y11zXZ9rhawgfs8JqWqpgglAYtX94XNFkKuv7ZesHnvzzySO3gfoLfdxeJh902CaXAFwp/G6v8gj
6cjvAYXcD6OsHTw2LmNZjVCDC77BE/B+EjefP+hOlUNc4y0MC0IWlEHtC8R/hwewr6nu+deCaTJr
n1YYCg/pd7+4YMNatlPZqcMx3Ox1aUvSug7uydeC5qHHmgMmCi3Kr8t75Ihy0jy+31Cw0kBJzzoK
f77yBWTSQuumc5M341CeoSvRa3jkYJqtXZOfDAlPf0u11TDZP0BADXDvkx4n+vddnRFEZZYFJg7E
6eVyjF3Sll9/ZFR9a5SxU+YVX6P5wYTPdmPRaL6EZtaNsFlK8GaSbNUhSVQHQawTwbwEihfTm+Jl
0DXE38kjmCWbddSIUhgMbbe61XhZ5LbbMmjSbieFKQ4daTZ6DPHy0WgOHNPA72qAsVLgm2cFZO5y
Hhzx0g8JA3GE14ol1Z+NGuBBiPL5Oqi0/8Qjx99Yc4fiiJ2U0082QYQTbge/aF/CQ3j8JeSqe1kk
IXG/b83l27AW6+UAykIUAssxkJYg74/bd9n4SeijYIbQ/tON8Oq9aGL3MpQXME1aIXnmqNpyovjE
cIJ8Ii0ZK894cB3bXOLdv6cAm3DUOfIOohKcHSyTejEUCW0C6HtCCCAVjfY9XyxjH9AMz9P7lbd5
Q5eBnS5jVWEDWGiuFwFfJ+joWnwxBzzOJKMMfdA8Cz6wYyi5oB1dDPApXmeClWMErG3AMCm4Xplj
moY5gjVgBB/UoUmtIboKcnqDgbopN/OZPEYyQil0ExXqkZWZXmAyWSNWvq3MUm5c1cRIKYX0gZBU
rzK1G5UT+Wrg/Uk4OtCEkTtWGnwnSvyKtBdIB7dzjUNSHq5VqKt5mm0KpJPfOyhzJ0AYJi9YObaC
lxIb8u1N8mLhWz7t0J3BxbgJBXAXAriJed+oEOz6l9c6CQe6yNeDjh789jRoQY9yXK1if58lZrGY
DCfi3rvEsypc/aPwgKzmrv71ujMJne7puU85ys73kKnG9Q7nN+uMQUl9EarJPyoYBRVjER8MJV8G
tVN9VYhaxDs0cTcxEiewQYw0UtK0fck6rU5iF/FMlzWu5sE/2wNagjhVOIJqDX3n01121Tkmmecw
vgLJkIKCt6tQMszgprTL/VhxwJco/URT3zvnzjXoUJ15KzjwFDI7xqvsYUyeHQkX3sxzmD5SyP82
flawh4TBArj5QrX0C6I80TDvP4YEInAQAp6RCApMRV8cMeNhHHv8BJt2rq/V3pJI6sfwzddi+UYQ
sVq/U8cZERx2BTZLiLXBjONQVKb0jGMGxB4l7oOP1kCpiSLKup30cRBjdJz6/Wnb8nrPUCx1Rg5i
nEtaSp6sTrbXYx8s5nbcBBx3WopKhxSz4yE2BqGRqhiu8Ap/maxJqYwzUXeoSPVg7zSDOyokrNRS
BW4LX8p0/KfSgagAwfe9aXP344FOoNzTCHjiz6pIGP/eXq5Upa4Zuiml5213UyK0UugUzy0ZWeHQ
NGHdqz0BCuYmo4eo/2CYBAE//7Le74sXVRSoBdH2E3G/msPNm1jq2qNaQ/bYOAg0ledu4OostuDn
syeOMqBKaQCpEpvvOjaM4RgGFNH1tdPs9G67Aq+d2CYPfx0JwsDWiXGTXkgUetoUQ0wtXPhvG/sh
9HJuZTBNIU4+XcGXdXuBq+WCZnkfr2KXlfEkYCWr0gllFlszU9hMyiF8nNKtDFF32nK3EXb2/If/
Kgt945UxF9ThGc+/hnufqRjBL2cm3wo7ehITEUc8Gouii9tjXKJlDUQyKO8LDKRIzDplJlZJLqrb
6wOzqVby6vijvOMxXwDi24a/ymtt7iEU93qRWhcy8m90cLm4vbakCPKLPlo2Zl7S4nq8gHVi5wul
L4zL1rW0rZvvoQIjWZm6rXLLMplYLiFZNxj0CPCx0sqomm8zryZK9l/g03ThzWOUG+gsnm7vFYrb
D8ggPnSCbnOUgRxhE20ladHiKBHd2yY6mJRBfZi37gdceUf3ZRNWOqush+6TiiOujEr4kvl50X+T
KF7RYNrMCAnxj9V6RcPZcL+7/Jclsnn0Tj09dsPrO+T5fHFF6S7AmfSNFus07Ek1fzXRMEHcKOEz
ubzwvMbFB+RIOIWks5nM2wbQ0dvhkQzQ/e0BeeyYVSrjl0aStMdx3sdpHUz/1Pn1/DnOk15ekePN
ziuyQluEmIeX/az5drBICrb8g/04mdQRvKf+EMpCdowZcRDDVm3jNil8t308X33eMZah2r8sWrSo
yfdOxOqgBPMlRzP8h//XhKmmfcfrdS1PKds3wGzb9Uvg5VPRZkHNzWfzeYbEvcXZD53yy+gnWKtf
gnSki3jrw9yVZCbGqadOzNgrsDptnAfuldwhVKrzd7uXsdMeojEOeRpSxNrBdxsqGqVu+z8N0TmK
gZVsmZprpCAejH00dVK+hTkr54kVIgUQb3Ilghz/Y7DwktHwUrFWlIUd6iBSC32mhgJYMUPHYQrs
I2qLAtQQByNYQRne7UVdloA6a3BkcU/ZkgOxFxKWfRfqXjmCt5l5Ac1K987dAE/LH4HYLUpjqUqD
zOyp6aTIgivF7UOFRDisZhyvBHIXydoJLWpFhh3ReE/Wc7MiRQ9M/W62fwKJqJ7vqILC3xHvGzon
meGVLoBk3/dDJnjgTrNAKA0WPEtcbAvA1Vo2rLHvWB7mJ25kipo6/qFWCa2EX0ouXRd+BAvk03BC
3YtJ4Lwp208Z82qjVFfyQqJZ20ZUGV+HR5dsCvbsbq6DMF1mdEuNBgUpwYKvONLwssku7tYhwn5Y
nPXktbKRtJliF7R7tKQQE2pns5XlSjjfPaQDnY/WQtfB+qcoVdUO2i5yYxjIHPAcNbyZInOXb0tu
/UvLiRnhnQHead+Eh7DLrty686L/tBSAZdVWqFv8YSF9+Hc3oXLu7fbnyAmluFkr9l7x6c04QVsZ
CZe94urjH47Lugar/qtDOF3TuYJxOzQhf09SxzZ/SUdBLNdLnuExIaiFpQMcFHXQbfbM8eIzP5iY
j0nzgkCxINvnfW+ZurwTvJlnc9bNY1qPGPMFGQarB3xFGOIYUwQ4XS/Ilvnc12GjYrwKxRR/Amib
mc4Q5q4ZE0d4V3uOwg+3dppRaU7gyOKiG77vUCWhaaWJAXBLjSq2Sl3VD6hZoEpYknA6ifTZ/Rio
h6Mn3as6PEMOqa3J5h53lVIExD2Ai0LfvTLn8M5Tar9Vo88aPYfRik2lGBMGZL/yZXG8EI8Qrvo4
2rY53eTVtAEZyZhd8F1JjP4/IjZp3ptPK0HuHa+Yz29obC4XWYbrRhfeu6GIPuUIDi36fsdAtcnB
YHBdHbpvuFWqYhfFCBtx47qlAI0aNxSmAWdllAc+yNYqesO4OsXt+w9NtGlesmR6AZ3od/MkBacc
TAe/Q1iH4I0Zph4NVxCizXw5ZSVdc51ZfiqJ3gnJgo6h2DRlvOC8U5M1c/JE6kav5MVUUE2TQHD/
QB8sRKLYhtsKLIvdErWUxse15QJXYtRKHbT7wNRT1dpT5wd8+Ad5q/3ipBOXTwpDRF+YD2XbuKhr
I/RqinuSeYVI/DyYs5lv4CZOLwD3MegtkZRKyD2sHSn70twgntTMQcffuQ53J9klfh2yR7PmHXVi
TsAE+MllFi238yEN86oSx/ZVvcPioWRpGnYyqMNg77TUK4FbpUeNpUF7gPhDEsOhXK4Sq855AZWs
+yEmMmQYzgq4gqA+trSLJ8fKeOKcAweQ91ZO8OCyelPGnq2uw43OkpE6c0slm7mD7FS0etynhDz0
j5egYyZMGWtJYs01OpfdKXnIFFsY82AzxBR028kNUBSpc67fufkm8DE4tuHETgceE7VwBsy1FuTk
17b162ZsuYt5nNwFTXefVDzhRQDQ+zEICIP4WAUr+003v0Uwm7Pl/KnQ9UXxfro+DVNEeOi9XOfm
W8LyCfubnTcxutxm5vqLd0IOeKAC50nrXeWzkHKEvrM3+uecSwGDsc9CqssarfGSe1hRbyXFFHcV
zBTPhSw2BZhs7d4/55HnBjirkOZG+1M8BjiWt+ZNkAfDybZo7L5s/od4Vtjsi+YvZ2lhGgBDNVHE
Y5ZfL7QYw0B8mEZOZeG88KFfrBNj2nvf4KJ+MJlZcr2to2uG7ZAm9U6f7EuFUEXbYiw149DikUiT
UcOyv2K/xKHAH/ulAmWoN6rm2JyOI9F3EjdZxJFzAqcBGQlp7FFdYgyBzK219CYXaCXte+GBljXH
O2UkkuYn9Dne8brLMh3Tfr8wi28a2HaP47zJIGdEqCZOsD0tiq4yTGze2zAOojwWyoVMwfRaIciI
Ewh7nTi0YT24tlsxDWs8x6N7hnQrilKvsdTInqUndumuNPqr/MjBOTclr+ooVcPLpb73FHsp7G/n
PWQflZpD9a1KsDAFzxgAeIugaxsgUbN0CCHt+eEGI8QhFDsNLFPyVwsa/suVVha6SjuOOxPkISN7
4Q9Xt1+Ig6HP3Wg3AvVoRERvOcmLFA05/1QBlb7luNHY6bianhscocvdxF8EfsSssvr379P9M6/I
hzsZOr0J7CMHeTIsactsKZbHHl2GZYPvqMZplJ0S8kNrDzLJMZ5OLlF3HwHhvVEClmiyIK8RnwZ3
1huO1DQwB+/lSMMJChGPYSSHRAYI6m7DEfj6rfE1vlgelnzzeM58AknNrzR+ymm4iktqMJya4Srp
S52s8PV/hkCjfsFKSqgIkue/ptU/HcjRf1hMyLBi6s4IP688QO1mFyuTRVC9Q8oldTUv3T/DAZQG
ZQWuES9aVI3k/mexCsxZp1oZ6YJG1d6FN+WnX5S4/E7IKE+o70zh5oXuATjECGi43TV0Dh2Pdpa7
OGEW9DEMgGQ4PTj5oh0AIVNPdZxF6Nv9GHMLYGh/ckkqeWfWVtxr8sVI2tABbkx72fFhrVp+Pa1M
FEBJu3chUomPyjWSnnknYRZbqjUUck5u6atI5M8YcCgpwiy8FkxsiY5lJ/RIdVwxk3Fs3UfsN7wZ
aCOQKuPqtEShWyw3f6HlFrhV4Hk5Rd9fhI8MW0cZtEacQwXXZ6S8YPx8z57So4qFW278/M2t6X7M
Kqt29gU8oNtzyuudP/vyHgNxDA296r/oZX80b3rsfHg+vG61sak+uG1IdXUeywrsCudud0HSGr5M
Mn0+aKbf5HXmnVnePhF0GgzPo1UO51hsFkCYoROWJdESFqdTl4zuYFEt5rppbl/Cxxy5H/sVLvYA
L9y7yyWB+kFl9vrDCJDzFOWnbD5zrcIxytgqTSNledAKNm5BEi+wv0KhS3wmeCrdQO7iDJ4NDqNT
lrcHFPfEwZuu5A0JgRYCoycQnk0pIBz9IX5WHSfcJF1s/fIE/pn3gtsroSiLNXQlmnCtXgO7pmHd
JQ6uuzxbt7LOIX4GrMVQfVwr18TqLJmouvTJ87bNoBp2s1SSrFXrBVJsHAx9czcfQbmPDS65UarO
aPb72x63dJ+ayyHoZ3XiCG2NZmEbNJadZmxoeprvgbtX60GDx8sK95gUUkeQsxcsBI+bMl6U7GDC
+9q8a/4tmZEdHj5uTTF8AgPwipkP5H/FWEIGfxUp4GQjiF6bXxG51eQ7SHrwvEzdFwOVRGjMIkJr
o+eeR5O/sUt4b+u5MFmvP9ZZrrlAF/DBtvRe2wC9qO+IntkDWadLIoBvmm/HibPrWx/YrI+Qe1fO
3VZ6nnPZymfDh0r+Ea7KhTwLKNGe2snQI5bdNQygzzxaMRUBc+n7BrK3hmVLzWkSGPADzzS71RM1
5XbDVl9bnPn2e6Y9Rz1DrBqsDMzlyOXW3K9xyVePBRTClKvTndFypQK2rkwnQJmqfMXbCgaCaIjB
b3LraZ+RAubUMhp3rTfTySgZFtO5qkN9LpmiZkt9p/urKtwHR40RkaGxxrF93LjtUtmYibYNlV9z
mYrvTtdKKM4Yekmf77lcUyFZ85ZGv0qMIajq+ahaoeYadoEm2cnZfnM+jnqPEkkMT5jN5B3L+otB
UGN2yFY8UoodZB5IPVsR1gKG1/BNOKEY9Del5pHkzLJgCZviXuiqcveUM0Dc0Lb8UvRewTw3QjFj
6kz6urFYYKsX2WSJwrr1uqmgDHaSCMW4WkjKyizJZKmk9eiKWPLpEVqSmflykYDOD4NIqEPZDWMd
AF7AnmrTSvzYoc2o+wx2HSwTjCb4p+ZVG19Fjrdccn9rzYcHNcXldOEUAHIYBcocAGT/hoBvHiBI
FefbIHlu40MFSn/WGFc6RYu/pYLTnnMdwaXVdYctXT0ct4+xVeHc296J3q7PT4bKFcAy9KKnAdji
CFgwSfHeNWJ5EcqFFZLaraKJ+9Hx4naN+aRrJj3cuB2M4mr37zoqqKFabcULmMMOlVp3KnILYznp
m/isfX+NALT2ZB1/TF+UVb/AKa+5456nvAhw37iKnCQvQjG0oEsOQBcz1tivn3PQADPttWqP4wqV
XuBTKODGqwGhVHnPKr4+t2OltoTtO0dHrHGNwRw9pAEgxL71yM8Y8jAKjXI8ikQzNdjmAKhOt2cu
gz9T8uiPJ/J0sjeKSfSo0N3/fzrxWhCjxa9D5PCBG9himDpkzi2LI1m3u+fVuj8yNS7okhIgfd+0
x4Po0s1gD4WaVtpYua9+s9c7kLsH3iSxvK4fVjmZ3JU135HZsmkv5OUt/KumgROK5DMnlDd+3FsH
SNYMRm+kAN6zLzyvxfOLA0qx50PAFf3Hcz3GkJ/Y1REsItrnpa9lUd5MBFGa4E1y3eYAbZ+NkgD/
Dn8EaNcSjNTCchSGZZc4+CR+PxdUy5X+aCpl4mjcqvbH3MrMoCWvTlPSSGnpr/w/JXepDgGfvwSo
rNFqRxXujQZjr9rXQATjrdMqPihJsk/3zCoEKM2EIOBvBH48RVtDSc/bRY73G75Po3H9H2Jn26ot
aoWwN/c1+HdGsd8i4HBXWM/G3yYnJPDpWKgBBBsGrnxsQA0k+hI0tFn7vX+cI+m2W8VoFSjzFrMV
MZyqRZmV6DqDV1euLRP0Q88Wr6gAA24NkpE9kLaaLLcIqQ6yHFcIv1Pa5wka1Ix8Cvkj7eMQ1eMn
cCngJdcKwHkIXyxRPV6CYvm++X4ws1AahD5dgRYi0Oe2ljiOVu4ne4J2cT24qTcsDA+ej1Jw8aWy
tAbXKnWI+PO+uz0G6TQvT+Fr2g65Lsoqc+a2QJ7o6ocU/2uXLqemsa3da7i91KmzM2NPa4PGbiWf
BvPuVPrlrYVLc4P2rUmKi15NNBfLtPo/POfJwkWgBPagsh6cQLV+k8cKK37Bi9fJWaeUVxwPBLGf
DS2RBbAPE9SaOi7iipQslmlM3z4te1uOjgWYQk21SEHaw05eq78R6+Za7CBse8Qlajtf9DSLfIOm
9pofUBOqWrrgcNsEQefrzLU8mcO7MZHJXyOG7vXcAUekdNG6zFTOKPlZgMiwgdBsr9a8tgxLcQMe
Mi5iwJHbvy52SEcj4Rf24rlQtY9++4h9AWKG1TmxkEl9bo8BSf/fwq2kHIx6xf4k+Aa+y/+yPg5l
jmLaPftJGSGQTG7zKac0tdC+CbFuvS8qPzBtcnQOsXF2OEpZiQvqd92tZ+eeqpOZ68dgWbWEAGNp
f7dU0T+0Wb7JGjIWgFzBTFSybqOJ86qfETfwZJyQvQ1pfPEgKq4tCARDnXKLJxEg7UFk6N6bCufb
7epeUy2+1Xq1YfsBdbN97mjpRx9sigXgnBcwC94vzV9BjQqZiZMzKvIjVdizyadN+PLu3lweJZ1Y
pRVinILXuU6PdvNbehjdlt92TOj+K6RQ1FmXAjugmeLw+Pwsb9X1/K0SBWZh6UQqSMk3GZpHjOCM
VNhkUMqUuJN8c4Ru1NRmjZqm619fB73ugzi3zLoUYqWSDi31oM46VIYoxqGpnt7U/f0eMlMVMBix
xBbSaonjcQ5K1Oo1sP/KL46oxm4gS9An0ofHR8cON2lm+KnvLXfp8QwlPjTAT3Ymz85PWpIkVbVz
aLIr9KN3D3JsVTi2GvbLOyjdsDF+jJaFLE8V6PzKUl4t5rsYbXDA5YpDDL91uxS22golA1WPOPD+
2Qbg+rKhoHlsSNC/g+1c7bDJyrZYXLWEvhgv9jKiL9QQSfQC1YiZqBgKBSc5YxAWd3Ej06gpx6tK
nWCdYe4q7HOg80u+BJ62nIr7x1+JruT/Ph6hTv8IqJfpSw005rPMJuxwgS+kOzOLMdb6aV1AqBTG
U7Ysss1AkdpN5/Pbj8Et5GJ+5O9RHYJZWhIcAldcLESKZTXOxt3gK23RFGwyzRuYXHD9K4PlTHCV
3M5mVL7v8qIo2fXWUe8XV1ooddBPQWX6/tLCQ0WCC4dbjX85XDWVwflULT0kIjxRXGJJlsjiLRuS
KPKQ81k7VJd5gwCVWU0dvD60Ek4BidRRQ5mXxY3m3VNhm5ZnmgWGL0fQWv2+GdP/jQ82j9YB5cxw
gMpdPdmucK1pntW0lE9h2pFcZzpNITfBGR2Qj07k7Czt5s8bl6sTe1hdtSGfjzJ/VqR71SBEFTEY
c8fYABWW290ghHjqLwDB+msbbqhHkd+3J9iFaW70Bshq03BwYeEzuVbhl9O+DpxuBP9xgY+qjiJY
HH+lDc9i+jOZjwlpSQmBOAEkHy6TF3m/s0S4wjknQYHlPoEvMJaT4o9E6TZkJzGK1aqShGIvanXA
TG3t8WHRmmFQ/WbNd3fTIb7cJJ7ehZw/wPvlRhKS8Tp8uePX5mtTcUfSLMOh/jC0d7MRnNn/4RN6
6bumfhL4hAs3bBVtDP+RBH2o7iBm3hUEo9cRav1Ryp6mxYP6n3I6X0T/WK7hTYcQeAogvAcJmIqW
8Llb08SUQ71iInYSRDA0gIC/GOHxq1LAwYCPfO59VLPXYxrBLIseFREhlxwUz4Gicdaaz2A1WQ5v
P+SJ2wbh0j+FrwF6wo5E4oKN2e5WyjfP3JznOLfBnpYy//KqyEDrPJKMzPaNH+TeTV23xeY2bjCR
Me0xMbwbohL6JfW+ZcCZM6bu4ksg8vXDlsjtpvQMyJHhBvInhHGrqowYtJw3R/4cDppTcvG+1L75
ZtXZ223407g2ARFjMsXSXTDc3K228RKxkLMGads8XRJckyvIbTyxGRb/jo4anhHDETEYscfbsRXZ
ViBywaNd2I7XJfvxJk6O2MEsfJi0Q8mK81dfElQoMzurUefqvoZXcCRpfDyCsXdd4AFvh88MLIdZ
A3rN0v6Ypb5JY2j465wfd6qSInhIR9EeFvGvhyORkuCX7DNy3DNuwyraqVFoSC+yOlz2bnYmm5vK
3ldDUVIOIcrYChsy2aB9EZAHc2LzjGUM9LEtX5Ga7qteeQ8Cu9dayg40FTSkPgfYzd+qJ8Z4HtRP
nvh/RZ2cGRFYvOAFcLdKTZyLkoZF/7EdcMiuGyhTX8f9DY0ooadHYwR47sbXZ2jwQ0njdcRyXrhR
71x+QdxhIg+SOqIFuzSwBgFYIx3KpvSyJhVPiK2qoCbboGUNZMcmRtTZvkv4aMsq/jZEk4up7ifg
UdhcNP8QFp974/RsK4iWum+PgsZkCMtT4F1DekmF9ReCz2MmjWkAtMCrmCr0lgunuhKWIh+OFOkQ
JpHs8fHssBesxcVDHM9YD7iD8Ae0baFKQ8uQgzMJsKTXpz+0gcJ/ykqMSJoe400wtUlGOmYLDdGO
2i/sxlezxIQe9lbqYJe0CIpzRZPm0Jqi0MElwl9y22RtzX8+UZE24MVqnzUCnvpnLxpJ8QQFii4b
qlaUmIvXVE08k0Kc+eWAYCAmrsN6amSEPt2FFQOD3LWI9SCvvMTP3V7KDeUCK+YgIgvaQp2NvGKz
zwsSDDSNaHieGgf20lxNkFPROV59Q2JcHolrxXZiAXAXzVlPxwSbSjPnPVlXhMw29qP25vmtPE1k
GUxzaT4NnD+93toTa5uGl3hcjBCOZMDZdJRxbpeE3MDeZ4WMgorypDzJWPPHuWMv12V8+bhgWBMC
JhUWyMZ+1DS+9+SX1nCk5qj/UHfFa0Yc0+mev6jxzK7fuG5WE0uTb25nytUufTlMqzHJKgNQIhId
ZZ3wQBiQsRpIIfJUkpVfLnpMcPNFId5IDTaKP29gAFYpiEHSryenNoy2nADY+fcVT2KKWBG2g9xm
vRRkPK1PjnxgQ23JtUy5HlW6sxYbw8FSegngRiFTPJdBg4XHrO92xON0GMjWGK8ZPxAdJRiRmDqL
RV1IsMyA9zVOYOkI+pPIRo8s8TWTH008c+iqK9qedybXlXcJLcHWTHOO2uZj+X6+N5maBE0I2YT6
XRigSMT0HypHvZMD5SpM8H7KmSGn6KRCCcwL36YiataonlENSAL3L+qcsoqLHRwWHQWlrOplOAfP
/jvjX7bHQvpUFdnAdFLqGUpIkV9RrWZes+Dn/EyXf610ES/8yACx90Gi8aMzULMOoUS10oRtRc7w
dTLVkH5XC15eLL1aDqMHd4GqizbVz+UM3NXa3M8/bwDf4vUPHj21EjFIkLYOtdCsNeZcJrrpO8GA
/LvxRYShCqUmb1Eqs0Vxi+G1tsAMbZC01M5ipJ1fcnubLf8tlmPWV0GXj7zUXhnQDGRJvxl61pei
Z/X1wpogICQoK37RYb9QQFVVGFhGU8vcTwyMcgAyB2eN0LD7B/Au0gp1Pam+zamDrFehp/EeUkR5
oh8seEJcBAtYK8TF+Yw6BM2U0Kdq7IyE1qHNcuyzcL4GVaNVzWGa7CmIqcxwwT0PwKr78oVI6FPu
3ntAEYd7xDvBvmFx2cv5JOdQ/tGNjxdf7iaEBRwrPIkS+JYwhDeWxHB6fOZW345KlM1iTBfT8wXB
YG3xBAryh03FQdFL2yF7xlzv3ab5APZtb7jqIUt6itgPkJGSS9RoXi+NyS0R/zZ8lFv9emhs5KEY
YYzTywR7ywykkOOfRJnS62yUlU0v9MNJ9dnamwt3ACzrEsgQzpUh5apCURhVOl3pD5RxIsddrN6N
5xTCVdf0/LGG24d27+43IWE2wbnF67XyL5o1Kc6nSFCK9zbUvCBJDlAuC/YpgzjY02qZbzaPQ6Qw
XkGdm2p7ikfgaJvGEdcc/Yys3GUw+RTpuoJ5FNELwWbmn5SkEKei3ds4FTqMzg2d1VXXT868OJie
C0RGLEbyUCuOKDwXKpqh5QaZgNDgSV/nA1upRLSBTWAwpmQPDLDSQc5X3EJcjAW8Cwwvs6zwazds
kn5fNErJhxi2fsjQl1jkf816hHH5zGszthpk0205SNgXAtf3fSYwCKUSZAAMHqJjMsvzHeWh4UOw
bZY/ou1cIka1q/RqhDB07bNhH0SLOD+ZfbUq5PrpesSL097flbD5Wxecgw9PUXKOP3JFj22jHt2c
Q7ePsY9pP2CC8WLcvhGWG9NiiZ1Ua9cxI9bQS6X08ikcv/I52loyXK70VlfaJx5T8AOdT12SLKHM
jWbOPSELf049YTdU7sf99GV25+mpoZRemmG9faTzfihiMNxQYu7xw97oV6HCBiJ0b/YAZFo//cMs
8/hlgEfKCkzrvtGsOlUsxxEj5/i69jdtlGOx8rX58Sjxc+o3+9vr9adjQGerIaoCk2ub0WwGYkHa
U88p0rFXCAx9+fGv1B2DUhlHKpF8mnbN1zDTSbt3Lli5hby9g5p9y1fjFQlHfllcQ/nWInY8E4yb
aQJk8kgdonMuUc1uvJ5VqnHmE+OTsLXyA0O4ssX9+D4UC1HBTmE6jGYljN57RuJc9SiKOaoNxB/Z
hZB80Hi1jUC2qNOoYt0MQmnYWZU7Avoe6Id1sbbk90Bc6rQVj/wOH0ry/VeuEKZMObybc3quyabT
kSZ1vitm7yKONgTdRX7HsGrDsgAvHVppxNEvnS3mI/L+ocxN/L3M+Q7lIpKBEFs7QtVAYnnsCS/6
84Kw+X9Qyi/UYFjiJSzXFW/3I74sJUPOwFWJ6Qd/+4f+WnU71EqoG6fIc0bN6HHLwsCcWU8QjK2e
8ws8iLN5/+H1kTLQKjM0RQhr1XgXZ1q7qyOtumAcvRK9WO1KsedPqGhfsBVLaxXuleuRlOTEY9rp
IJ+bwuXllubFnBmyQSC9ghGuaacLdNc8+YiCQHXAmUlYXSRMCPrOC6lPyhWr4lyrvL5O7FuzqgC6
nBj2ssAbQYKvDdGRAgN7cNJu8q++avW8emubnywQPvzMbCK4zvHIt9ZClE0ZuCHmyRNedR4gr10P
9UKMs4UzNPIrkmeKxLDlnj5WQO2/vHde9cKyb2DnZq93YpF1gARFQbn1/4bMbre1405guWTYD0xK
dyoZdgZiyhpGzRLTsB7wlcb/NaCOMnYyabRdZnH5TRduDkY6bF2Cx7zlRWx38AUCeoOiQLFI4wKM
oWGwzpn//GUHNBenjgxsvx0j/7NPpuu8f4irdrkwCP9pJ8VFXc7n21lHoy83VAKRa5DyI/Z3EL5K
fLnfH8EKSOO0R+C1LLvQsmCBB9P4Z8DHJbaJbeJEcmu+Y0LOl0LEoln23Z9n5rmgvtY4aMzJC9q6
5sxOgodBdqfzilcSEj5Qf2QO7dKSu2GpCfshJs+eSxjPYMZC/oLTsMOcvqx2GXiSbVtnS2evLk9F
okh2H+9/3568gcyQk3jB+9R3Fv0n/waiq0jKv2DPzqzcKkOfjFMm7hZcb1Rm9PM5BGkxGKBv5pSG
R+Xq33MjEKsWy8r8jj6LdgEhPgWPcbcmVBeEMcwXqv9Lhl8GuZLJwEOe+IiiHL9e0sJDfh6SmgOu
3LxD0DlmgiBYytQcYVPCfKpDw7BwI6Zarq8oD7/MHoTvBW/lI8rYmv5PkJFio7z6wiDAddWO0Bm5
wwkhXqjThlT8nClW1X7E54wjzJzCKZRhaSw5VLsBYn71mSmSzetn8798NO6H4kdtnygKjo26Mj5l
WC9TjDVP3yaAJn1oZcL6x7gkNOBu35DHolFVmlAH/1Be8SZei5ARR7uKISA4KYOUF/owankakNpv
/jsunsNjJpvXHQhqvU/dXevpZpX64VQaQ3H+96rAC/nXQ0U0y80VrB4PSYvFpvcss+xsy8+CtpPt
QQoDnfkT1wQEEYYVZIHN3copi43po4NWeOPmDRm8GFBnUvvQaFkT1s0SJ8Xupn5yh4BkpuD9GCF3
+ii//Bi6fQ2COUrmlLpw+vuj5dHVYHqU1eOv/PKuL7HLCg26hhvA1TV3VYVapLqEBeXiS/s/MA+6
g4ztEVLflEbrmDjnwPDDhC/mfLi43zG8P1F45se4rOfRj5+Zi8P9t9Bu2mfQhQj19BL4CPryIikt
98S2XeDnAW/+m+SWdyCx/bbnPrdzWBFXESuXCYhHnyTEHvl54150NWIuk0S04+oa2BhNWu8tZox/
rhosWvqkaDGxKEFFQFY+gFyHExozghGBkKGYSzPoo3hZhXsmaJj4tFjlXIUlqcLxAzncOYjAtaPI
lysPMgMj9LL7+AUZskxK64AaebXGd2CSV5gzz8eOtTXsb0xNs0nwrmj5OB9RyK9itAvcfr+MhI5I
p9q7BfGecGf+IjIinPBxDpK7JoeItyBUUbkHmZGtXVmkPo1/e+6eDncDA/qDGazGo/v/ZbluuAGO
LhKQVnQ3IFLIlC42Qw0pOCZenbpS2FUnkMatReL2OUexp2D7kQ1i/G3Gdgl1nUVMas/M7bPrYi8l
Dtux57GaKpWrMw91J/nyBOPYB/sZe5fWXfWmsm2fJ2MCS7EPBTHGkx34Jc7va+Ieyi1AnxZ3gghA
O93veweoUXHuD6lcqpxnQgeX8LiiqE6GtT5G+dnPLrcpChduhR9WEV8pC2tCt1VwSWFYVQy3cmCo
0CB+yTqwQ9L/lVdAQLVTSqhzGbVxHnrlOm0+u4ReUXK813Gj+u+UyF8/IDU8VBVobRP98CKeVCCi
XVfcK/ypIW7a6M9FsiQqnUKQXPsxgmLhCreS/cMdTcWKqJHCGUnZjgaPz7eTEakGLZEx0d/vjy58
3eND9QvXjcdu5nN0jSQJ6b3Cs8WS8Db4p4IZFF1Z/puO8nB4Q5YaQi2wyNldRH5sFKxNm2uufhHU
2ZD9VKV7f3QoAZmn8y7vV+ChmoCag3ACz2y0uCwDDJGq+jo7vXT9KQrUsu+gx18MozuoIUvAt/ZC
H4XerCIH+iTr/6eyhNNBjZ1ZoWRi1ARD91XVBITiGakDMCVh4Rj1VjfNYUXBXGq4NJQQ4odACcO+
j2WMgkC/kAHoQbUpQak4Ei5RYux23K6BlRonM2PCgo5WqrCsF79UhQQz+juU+APtyUvXny6dwkFQ
VM02NdilxlmnHBtn/bfgl+N7Gl8X+knHL/aBr0gS1k6PtsUYbOQY6TAuP5iRq+0vLUfbbSh8Rbj/
jUCt+ZH7Pzcmmd5g3Ue1LSdmMNQ0McghVxOJAmvjejMus4F+a8AvSYfluyE9joB2In6gVvzfQBtW
VtZxQ1iDMo0tyUSl9oyzSIk16fgiFaRGp4QGHFG2P0Q8lSoAcBqOf0SP3AOPtJ3frhCSvj1BNAQe
gepQ4jiQblVy4xentkjWAatUQWT185+MTafJ0uADl0DGVC0I5MpqhC2ylYXIvHbvBNi0BXftesug
MOtI00Dm+UqnsNeRc1XyHy/C4Y/FJWgI+09UmNlUGQCpPWd618VW6jCecSGmBpn2pkG3qhHLHb7h
j8a8jST48RnNX8bnJp+KP40YzN9tO0ukTWRF5vTjTH0gUDI1CsKEhGdwXwH4FiAK7eBttmFDvXOP
MNYUUWA/+OuXPVzXm/6Wtsji+VGQ1J1FEfPEbk9qHkH18rZiUnWRcDsz/VPpSbVl1wWQyZvjag7r
dnrJsRIrUdjjvwqUviUFQFRTtx1dVZfmMiwD8exNHI4CT6H8lz89WydkveuXUFnI7S0KIf8F94Yi
faoGrFhB/7IXybMC8M/Ue2OyeR1NLoFNYzbeds5wjRf4C5uUpxYsKpXuBS+nxypddsE/EmW9zFa1
svIuDfCzSTBGIWyToRMMmyylVSxfzZTZgzb20kPczC0SbCIq3yhUVJ4nZadiO1e1SsoW5Mp0UBrO
U4SxD+PVMCNPpHSnjy/3c7d838axUgtwGpnp0gIOxe17zByrHQLfvxOpSs3ZnHn7LoetSYvt6lR2
kC3Lrq0gFtQwCn3zxZVIFwwhx02XYTyPI8Iv0oZPli67tfdvAdyDmooYUO13Fsfge4oYMmdGx4E2
FaZNv3ez3ZvTNCyxA06rfnBR1bkow/5q+g40ka3T5DN8Qtlpr4qtirhdUPKxoZyf0aPpywWYfKwK
GlEZ8YpDeC/sDQvLgSX2Mc4sLlliVUpSCN/+cRD0BsnIL9xhueNtUhSKHwQkCJP1tOliv8Vk3mk/
uQtPPhtP9jxxLxzI5htCbxATglqNLIJGtgihBj5hMa5MZkGIiPNBxp2VKPuj3AIypFnqrEYkbiDk
UfCGcoMypX0nXE4mQIeCqxrNgOkSqGXonxT+/arW2mjcWjssuIYHIUyKols3FxkaB5uN040hettl
7rHgaB1eenfI3xFNauIGJH0R8GoNGE5PYdBOC53nLCoZ+tSK5qgpTLBWtZxkZk5Pa1sQ00qqAO79
AmAGxowrbdKAONicRTgI4i0C/JJgUJ2ks1TJ7m+JNBsfTvUhiPIaQtUNDyq1XJpSqcrZdkftbrSF
P+Gz5NQsUrFUBkPztmUiSRjHL7jZqaMomgdBzCeP6uxwG6hn1sjhUl101s6A+/0YQJi6LoG1l1gU
+rbw6ZlkPgo38pheiSSQCebvdoCmrooYe8yfklAA1ECfmbWmPPBbyaKwF2q9VL8KAQXFBWwx+/M+
9oqKbB5vbIiQ70Nx0kWbemV94U5RJf/rkFLH5PF8XKQvB7hQEWqYY/IKIfhaeJSJmbKxxxTsKg3d
tyjcrV/pFHm8unnazuvrw1VNs+ci0wV2HPDN+KaShbks+LoIHtVGivaF1M0io6OL8FScZ34shNwS
MvnjtQZbQU0ymXNw1v28i/VTcDC0eNEDReENFFFW7gOV5ZmKksUaR5f1gAs5GGIJ6fCjIo3UKYJa
gPYs3QbOY35XqvL+hwqNnyyH6KkgGJgk+/qTb2p0EOzxLeWdXB2E9rGRfpLCQKfmzgaNALcvNgzw
TfSzkwJ4usQiE33iblyUV3cnaoK0jaN2i7R90VwJxAxASPGMethdKFrxcOxGN0qXXzgJoYhe/+pG
3Ycq2hubmlcnPpVtTpRYdsusoXTxkGbj7g6nZyaHQFyfLvkgsVm28g6gxo+6jPyTmZ8FDNFvIfZ+
Pt2wwVrxENIvGn0njg9Pugi7s9ZlQK9XVVia4AKQiai23H7h6wfstJMDxqvmtsd6NrRhey/Z1LRK
7ScMPFjnhZvDeBzrY+gza4RkDXMhRfIAijxS9HL+Hvyec1h+kthJFwbMwhLFupgS4c+pLRFRoT+L
5R7/8xYrBDEJ6hR+HoVF49vYy251DFOefC0dZpIhsXBgn9kiqe6l/DQccDTFuG+VvK3fhOiM8awf
QFSH0GfxP0kRCBeMux6+hc0csPUCyb4RYNEUU1SiTjG/FqIk3q9xaedYs8JnhbAEvDN6AMmdtfJ3
rSfWKxaSOgnZuuqEuGw12r8YmAKdow4hni8SlNko0vScnIdTnlEeNtHPjYoXRsCg2b2rXzG1vS4t
KAdJr2oiI3SIIzGL65rRmZSBhA72sCRcpTmz80h2NkjLNhp1TVU6wVWzrA5Vh7RWzuvi8a93hXpo
cu3HmxMuLJry+OlzR8Dkk1MA4AJpoY5GtLdl2YBIJ5AWn8i7b6AeiZ+5RtIfce7+muHl6IrYO+PI
Io6FOI0LIkSwWZ7nGjrWODG/GwStf6qLAnOUDHmtyZiqvnisYSuXsQYlVoNDVnjq1XwawKTKRXF9
q+lDLW7xl54RSYlw4RZYb3u4JB4ulKamZQMNYVu0eiQFLeDaBWnA8LfNcolTEKqB8hTDyIkpiGG+
UGgahnCePKXaGgzkewdwfC2Vxv96x1QqrryjaHCItzsC2gQrX9GHWhc8uReNcJakw8UcxjnvHtEU
wgp99tQD8PmstgqDInK6SiDlteal0+BK23jlUmG5Ibr3Ax2ztT1wAM2tR1AJJvCqgmV9N2XD+i3t
Kkby7uhw2m8WgP0U+3tf0E7ojn6WjgZtDlscTFrjJvPeUbEmZ6H8jBcNhOo9XCnqc50nkVEDAAR3
Q8ThcVBnNUrLFji1jjn1Z8dwHQqG9HRz0PXirvc9pFpKkf0Fj8mLuE9i0GxxfanGSRpcZN+WbRas
BpdN90JGWxsWo07oe6xVgLu2Ibg9HLapqiDMdojx3YHOTyeRlUD0wCLsrstCliRgQRnlWZtnH7UA
K8sdnLiKcETiiTm0xHm7EDqZNlk3/CWmknJbREyk1mvLXYQursniqFA+aMW+23Yr126ssREHCWyP
bovFefr3I+mDH9CzfNBXSVRqHheNho8Th+tEwvQLKC0tceotlsuQoAxj43q7iJjem+BmEfXytLrJ
Xvk28poQv/UHWFtaR8SOPaxoUHfoA2Yb6lj8guGzddPJeEHB26250kGr91g8gc0ACATu8yTTpIIS
DFlNWNX9GbS4yxNTBnmPb6EFBKBBiAoW/P7C7CY/rzJ16Z2stIOScJsdOeybfEmiaLUsTn/h7CMQ
uqS+6SiWXhvn281mU4qgF9gGb7uT2gBK/U8wsXf81fv9RQFJtg7CTdQqjdnLrwUAqW36CkDas3Bz
3trVlLTBvMvfRADNU3NB/ft+WIymf2y+H+bRK0e8aPW8W2vH1ARi95TIRU5qRn2ySGfvhaTAL59g
mJ/Jf9q46Z5gPm4ewl7f7mbScQqgVZqFFWCCZQfnAAPNaTsdSgEJLMkhxfuFKxVvqJdA7o2oDb6V
RyuNM5LiPSNgf+uJqNf9RU0fLCFm2YDrmLPXZDbPOYW7nrIMjCRxy9DX7wudlvpgsaf9i33YyqPh
Vhh1e93NJpqG3yBs6VS3XFALR+hWz8AoBVENSIZan+tYzW2BVeNuQO9YtqPocO9yZW3jEbs6jrUS
nHE5se5g1MKU2dpmH9jPkusXjdDGyY8g1tSdI359tW+tDiKqhswcj+nGcJ8qgoPkJBXhOx5zgYg/
qApjZDrjT/w0ltgv7Yu7hHiEEAYviTlFr6+CSa4jJDtSm+o7YTFbVLrloCRjwHMs7N1+dxY4KSRl
zC+l4SutKnuTiKhDfEzasM6tXynDdwz3FnYqefRwTWwEgjCmL2PBe0fpOUu6dTOn5K567Z/bm5zF
T+6jO2qmJy6t9hswYvYi9Abk5W7Q1ASvhH71vSdF0mbpbCPc00lhLKk0cbJRlZWaGJH9MXE6U3Bh
6sqPXaxqTy2wyxbzc2mjbUFA7grPMLQzBFHGyaWDUyRTlsU61bI2uQZLYvpcyG7Kwi/JDxMVL2U1
CZdYA4TKSjkBYOCOCScelo+OI98TN+wt6el0nha/uP0M/JAjEWnG28TxDT9+daSMb7JFp6RGzo0f
rvtNxRzedPtQbHffscnbEL9TfVJYohsJHlhDGbFe/5fiTKo+G3h2kW5ZgJgNuRz37K8GY4azZNnE
hP2dehLa4sZcYPJ31/qCNY5YSBFVuoclWAOgVoOefcA+fbH3Uohfui6PfNEUWyMIvat5cM7pNcP3
rAH+rMrfo1YaeBCsUXQU8GLLK1eqqwDhzcLQ9yK3DhNyyjOsLsUMjjOUGsdgylTWH2zlTSNr3oGT
XX1rVjWZt4xaxFPqVsGRnZdr1TMlPYLI97TppdtoH8It0UHeFANOF3q2XLK+A7dg0yzQkvHerB8T
K9loLBrF4HdAM+lvI3p9LedrhVy9Rdp/CXSuHFzfyYAWY92kr/joQMqOGkfHkQqXWtWaYRf3VKS0
Pnm3l5KS5wczG9WaIokOS+bTO6YFqbc91uW+kzvKOyfjEbnE/O/Px+gNyoJgg4u2PhaT9BzzxfC1
Cjt2/DsF4PCGwKdKMCPeyPuu3DzB1iRoMbVYcwgpqo5NHaTCEY1XnhMUPJV0zOvA/QeaWaarfd0Y
HFQX99poOQftQm3mnz1va7ODx+9YAHaSaDCA8vg6Sn0Koa3vNgtmvJTXMNNj2MP0UnumKn4soHPL
geSySDcsUy7NOcSoksNqnTEwkH5U3JovQ/CzEzThjS65mWi4r/tlydUvQyH23PS3M0eQLfdH/g46
NbrLnDnSbyVhMcfa2yY/2AKFbtorxS2wuhIU+WwH+EzmNNFkCXEUEeYNsp4BSoJZIK0PtnathouK
OqhebG/WcA6a6leBLWr7hFRc5n550lAPGRISXg/gRhIz6GZoGWB+LUEyoxXv5DZyxjVUlGOe+Rki
nga1HFg14oSd45FAQgm6RjBvSVkc5LsLjATvRe9stY/uJrG73xTkg4COBeXqg0LEzijlHOn+Wps/
GcZxH6L542mLSJ/7JGLpoHityAeYV83jRQqiAx1sSlK53qzhbPvN4B3vcDv4iwoLZ/cJYACIq1EP
0014rEBc5Df4tmv2ba0d2T9Tjn0Ix2koad5g4lrNQg+uv/L3qM+d3aSffccL4o7L+8r+mnuaVbgA
vNu9EPc1nl0pmFbNOGke4aoSXkbdfNtlUqxnvTE8RrD1PXbuEM3Tmg+wVBK2X8+ZbpxMyVGyV4BT
ukSOaIj/VSTNNo30Us/lyYP3dgIshmyr9/DdTzcGesZJjR68TVGwkmjMI0RvBlbSRR2wpZ0aMA0u
Mowvsip6p2Omo6DLMo4WJOAB4zyStSjKIGU7xlrF52gz84on85nA3wwwiv9ihLJm2S0OKzbwnLEs
1ckckuONr2hSO/jUJZLIrCk/PID6LQ7961vVFyhf44cKwCfienxLgz1fLk+9EnEeZZBU9/QaJGRL
2wEGRl7J5jMfWCFx+kc21b781wZ6aX0J49cHyz4SsUbek1+SkeU6+/DQfJfHpOXVr+qvv/XXUTRY
n2nfEEKbV8u/rFWsvBsSJrNyvPkOV5AhFR5M3x8wbzdx9z3wZDtxpY2yDfRQ+U3Ha/cqRSx1nYAZ
1/gwKYoN+DkwQ0+3b+B28c5kLG/cTjVeHP3ERCorxyIyq/aDYaJOcZUjo1AxDKG/UX9aYF+9KvdG
1PHP+yhmpMkaKicZVzYZbaB47FPxY8Q8EyanagibrgLOkGuqhsyZnjxJl8iERPlXMCCMgJTJcrhr
wNt1ZGa+qmduXXpgQqCHa6yLrI/r9OUkjanszP4TRMrzveJjT/ZeXaMD7GjMv3r8ywaeRq6KHLvj
VWfsmgFa1S2zQnfQQCsBsT/dH6UM+w6xcIfGkfc5BMg5QBpvf3YEmK2pF0oKHoc58ezaTHOXdIWS
+e69s77qceIMZZeywwuHkLo2RIb1UaVicDisjeD1RVk/la8axHkIHa7cq/S3uLPJgTNtCMKhELfL
UXURkSQfWtO7Q74QKbfokIBx7lRvh1zhrOKMnclTTeWBRP/23dxvu7hID8miRH9igZy8jdVuWF4d
eC+uI+Vv29LLrFyY9Es8TkPNrnUPRxrbjvFCfLXyeshFQONZFeifvzKnyj0gIV5hBYxVAt2GJVZF
CK98j65xl6tdJblTMSTqRAcy4QfIZ5zIV6NV8NDp7QpTEJt7vVJpz++BdgoJDFQV/GiSvFl5PsUs
ppaICojVIbx2p/t9Q8GMV3xPKOVsPP9+hJA7pTIyi91Y+xCn+wafzzxtzgGeJO1nUSVcc9iYcKfC
HNMDBiMbamcLhgkxmf/vLhwOLehpzxB9FzndX9a3prTeYGGcoJBRowrQ/EJ+hijjVL6Eu2OS5eqZ
wzZpsrG4aXzl8/A6xQ36DWqwacbJuJIcmMl9Xy98Ag0OJAcPh8r+5CHDoFQVwPR2V2o14Q9iCWXd
2hS1dxDGTu8XRubmbrlzg6m5PzPEaH+CMqfZyTW8IWNy6AmgaBYpqdf1wcMHFbzlmHaeC1Afg6hA
00CP8T6EbtnaMHa6MyN/mjQtmEZvcRVuPf01cudGL4mmJymUFcAyoZFrTRWDFGeZBs1xulb+8jVY
f5r/xHx1RjWFPbP2zy9rYqPoSY0WA5sr6nxLo6hJl3Rpk4+VBY3yN0l89B6OvAuPRbH5hIv6YND0
jO+98E0be9QjcGst0UvMMROP6QWrrWv4HWBA1WVuhotb7BZkeLjeKEQeh64PECw/a/FWAjWv4m4H
bTF+W5XClUsi/ZUBY4xgIhAbKLStGZlhjSl2JgQ+Wfa2btGSsYCUwfGMFLN9sguGYEM5nySqiI0K
JvwSzusAK7+85N0ufYsGFP9cyntI4bONUGKOLzfuf9UtHkV0sGc6b38/gzQcNri2TROLcK9I7uIM
+fPkRMrQdwG1IZG8baUEM/KVbQd39saBfvAYMtayvcJQJzDaXJpin56jy4N24q21naWxcwvielHJ
uuFDBx22+aFB3qYvW3BrtgQmPVTHVDG+eu1btliWR/nDbMfjUDfNK+HDchTHyEQdZ04W9w9CcEJq
iP42ai6m4hu2g21MnT1zZA3ecdZ3t+qp83Z48l8Mxts2C8qZZfL4IHCb7aHN3+DzeejBVrap3PNz
2BEVmMFOLqBK6FhVs1tH2J6TKlGgu5RD4yJGrrksm+BHohVLFiIqI+Y3iMKESkGFJgJ89FRwGDrA
PNhhrkVC1oBoYChVDJYNF8rfPF3TZXB9nPFhKgp5J3aaeVDGyY+vNzEnqisWsgrlyaBOftgk1Qgn
VXx6d1Vy3v5VdIq/RJNUpnTXRZH5ui6fzL7f7yh1Ge333dtIreV+p72hsxZ763sPQmola22AFfXf
7nkehaMKs3thzlILsTQnIi8cMglWGfI0WhSC8RiZOjBQmFSfHhpiy8qwhOCciu3FlpGuy6QhoPxK
zmR3gwVhZFGQkYbB0n0J02oHnC0OIOVfZzFSRg6C6fgkVKXqhyRsq7nb/1GfhhaZgteqWx7l0q0x
UZP0OORXwJj0s+Nc+KxIojVb2JAbi0ZRjp6O/gdLGCiefKHPS5+Jg3PgC37QYN5u22qcUZPw9lDB
bI+KXSEdcFWk1R8VS08MCr0OVQ83OwqarpdD4uXXjn+5CBpjbIR4HCZOg1+GLvCqap2jIP6fcEZg
ZJFO+3UtFkkKdntoTBHVd2MB/8GeWteeHyly37uD7Nd043MXcLvHrQUpIN+cphvmoq1Z8F653sFN
QEexLh38m4G8coSCFsYUkY+bk9T2iUN5C4hVC83hv8a5Eq7c+B1UUy0VZom4JwsgRWUGsDjv2DcA
3CrrVPVm/LXmsnh+deC9YdKz5Q/eaVPa1z6hPwC2ZhsjVHzkTmYmUiTaXuLcNOXMEleY5lDqUuiL
KFxrnFgAk9eNKVgO3rBg57nt9yDyM+OIKo4iJobAQLAvtzviAuGMlraFAhBkT6DB8F1U6N5y3qFv
0DxZwusm2jEsYy58XsBwdKEakn7ZfK4Tc5uRz0EwPoNPPJgUXWiVbDEQVIhK2inu9gOyWzWVZs59
v8aQ6+TelcKQtLidkBY/5YEv9/S8lpiensFbH3CUp/uawPy7Av+qKfxZgfdsGTDopmOobqY13+mO
0IouO7quo/D+xtMiPaURVrlxYu1P/l7/lJq8BJkLxXHt5oW65NSajwLxQKV6nVkKH0KzpP7Ci+61
65fp0mfL03VHxsv2LKuaQkuD1/hxrClGUzHzEmjSHaUg4cTo+OY1Yu8SDEO57EWipE1IsBlyLKBc
ra6LNmp2D71bWMInqVmhrH/BjVhQX0pugTnYX37fJ52PQ1Rx7HlzNZWrtVuFr4dCcuorGIc9Bpnr
wjQiOQl73MndRhUp3/OeFfIvCmxDoGDAX0wp9oq3j459BDDbaNwzuOsDLdQuzdfx0v94Nk26Ib28
YyCR+KCIvenJ7Dwe4LEwy3G4Zk7LbTSjtF7HGB5tq6mgxBKrGi1rlURgJoDB5FVGF9iibj2Qax32
cbE08eg4HzV93NKMsMAKTIrvvqI/NfBuROVL8/vXyyIROIUZMKq/a8paKfZb/YdqwSl47SWNdEFQ
l7jcSlADo/eG+GgfrDRoLkFdH7Anbudo0w4lLxULkL7BaHe4WqUER1N7r/sIkDKwHETIIaZeeHcp
DJtESX2cddKINfMqrqV4a9z/GrcAPxAeWMPX82h2+3ELFbhlVX9Oa/iEnoKKAq8VsBfgjM8ykxnp
PQRQqsRFV8wuQnY+5IOqBu3E1SbodY1wtZawO4X22Q0OIaD5PHxlR0w0+f8SdJeihpTy+KlYU6WX
XII0EifoVtyYj2J5oFginQe0+PJlzecxRU4XTukwphwSjc2B0GJytYdf8ReqKoQV8JOVTA9bCrKK
/K27HlpRqu7QMHSOQIYrRDSct4ylsuisoNzk+r1klxhVGxucXEXDOdBFDNUvFfw4j9XaUzpg7ZLG
V25CmsP3LUvA7pisjM9yAuyKHDzafysathqw3KDnQxsEFXHPqZwXlAJ8mBQQSvuJGfacOpTXggAe
OaVn7wuvOGvgIjdyu+9L2AGYscRXvdwhOXCl0LW7xc3B9RLUmdlAbS2fVeB2kzfGErteZ9d5MUvE
KJ2I5TH1+UtcwL+yiGVyJOd3p1g2xD9ewEA4D039842/c4K3ZajiZ2VIMelb0dTeewPDDeiCn8RE
vher270G6megUd4/xSz57EH50wZ9gc0VZGgsY8AvBn9oZ0jFkreWsNQ3jf/0n5DuyhaCt6mYvpdf
fYqrdiKXDryC8+ypa1xm5ZpXhcPYes1pB0SXCWAQq/858uPvNJ4CYmH9PRhrzX5fpljGFvwnzpxE
ZLN12CbVd4nPxVixk6lfN9+C00MQ8zloa+Qb+i4ORmUbSP70k90yJJOHffI7DDAyqBjO6SuCn9Jk
MMVPgt3d0pqI1bVkDKxmEk9DLdLF3zJj9zJ2/9qJTxdfFH7LLG9Icwsgtv8sAn95HmT6jhuQxjcC
VcCMuNCchzUCOZb4VdRJCZEOQBmjZ0C48D6UcJTNm/+KxVjd7Q/3lhSMetvNXBftPnUE6PaBuTpf
eyucdWlOsVknGnABX9omDuiitts3mfCp9PwqI9cWJH/l5+x3O1RxQ3fCYVGi0scHOozLXpe4FlJT
i17oCT+rqT6o1LvawW+OVUmqB+i+omJxzKrchm2rBsDN7u+p4NF2fwrgGet7N2OW8kpOLlerH4Ia
bD2b9cKNk4a7GFalNJLQFVB6b20s6sLO/f/I4zd9NOP4AJxoMSlfDSOSiWKtlta9VD6GXhhvsrtv
0VFurnkCN/bllhB7g9oK0JUrXThVB/qY7TYBfCA0yg+/0v4joMmdTrqJIWnMqdgsPZLg2dOVRHA2
vPfngIhJ+AsokBG1ajJGzVmbr24rdAhb0f0k7p5nEvWtIgemCvcMabOCxB8wobPFC51uP4mILnCG
Bfy8T00V5oe+LkmxuJL04QOKSwLDOl7TKnZ+o4g8cPM++bpGoNqGBQJo8Z3fMFoQgM9YBhrh3Aws
CyaPeBEl7wqkiVGk88AA34p+GMHEyjbcVVPpJgxL1Q+150Pa41DWjmIyjmdwjq+ZAlGsApgrDKRI
s7dCC1z+Kk6SbwtOeY8f2pmOffXBFmzq4pV9vyHVnP0+MpYdiOEr3Uh4h8OJthmuFmbKwkGAviaS
uaU82bPskEpNOaaDqGe8L2m0cO6seMlgTglubqb/5CU7oICdnbdmGdRUYAa4UEgTCQ1pv+dKlb1u
8+uA5hgKuXyRDWkpdjtrpeYcgQfKaQc8L6WqS7ZjLvNpnkMfD7GCZQohgtwIxuU4V2EwlJoQytVI
SsZqkKvBl25Zg2VAFScpiZ+gtNoRBMxP3iAkdtkwwtifxlFveWD0nTMns9MKfeufxTJvNaBbInV6
Xg2NS+wDE0e2ZqDz8kTReMLDrAi7EhM6C22v0uCyBfwHA9fRmJ8OA73smMBDbv9naOksp4gDLOV6
jaDrhGAjEV+X0XdToGqd9QC82zRqHoSkAt2rxFHxtj/0kxqsdvv8b+YwpWgLkBnXVhQ07ilbONW1
L02IUQsSAHe/rVOJptYOlOlsL4tHG8dMaHLDkBnOJwCVBkLV0AwafiGdw51vSrv80hbCcEVKweXq
YLCbbFcqf6HGup82myy7Nje+SdEZ+QMBVuii7OfCrT7OOfCAFY9qZnlVKZZlutcq3voggriARHsy
xn1bYckCGDSaHgsHMLELF9POXnWbjUHVqpJDjKQV7suJpeD9TnucB13rG6hwl5uiextAuvn9G4PR
12O2IVI+U9rD/Xtwt6/IWcFHQ/SyHbGojkH9R6rvuLcwJB7JBtxts20wvF5r1K/+9XQ8nWji9fzw
QJQZLhJ96I9qpeb3LqxNwf1snrkX2H+eVJJfZSqBfCCdXMUN4JzfLQYF3BY2iFUDs3Oe6TGVgqkn
haGkQ+WP1YuJwwMx6RpQdWaFz+MI3721cWOf9rATvTBQwkXAGXoD8LEaJSgSJ65nAs4kyeC+3biu
JxfAD+U6Fcz/Mo/ZcSkDYglYOWqisyYY5FTJMaH7GzkMovWCuEtDzNt5KvsI++QrALuX9kzSYlN2
RZGgMFzisi/ESyHo3TWWtOvV/nQHAYdEqGRA41ToHQIhcNcK1vAbR8XkviCTopiQreeAoqJPl8gx
vpKG/EU49Glt+8y6103RoEpzL/lY2/bEMArrCWoO0WE0S2LZoP/3GhZCK/nZipkwgt/6okTwnqXX
jcFXojR5aUR0ptvCdaAl0JAhQy+zm3iVbJhrI+nh7/F6xY1j/L7zR3uIWgymAbG2dScV/R1CkG4K
afqTGIzYpjFutakWVbYOG7rAoqYLSm+mLSLsvzk9HySTGBENqbdP0miqta43jFON6C9PpqVqgG/F
6kHbgQN2leqGMDYWRtFR8E2Pz79e5VgKIf+0cAA/yrU07fJrMm5kOClUb1PtB5+VgDVyEG+rqRSE
vM6pSzr5Jkoa2s5TypOFzi1gEsLujTNBY1M7Tab2lPmM2ktBgqQIitseuVZMFn/9o4f1vIyt8Inc
coMnQEnqMMlRh8gUjquKRLGZj3DZlWwfrE147y+dqStuzfxN0RHHJk8BllrA2dmj42iK4fkkvUXy
1eAg7D/mmZ4QKjvGprfI3Tqe+sSKt3nBtK/73flPKss0gNa5EFv8KXXkkCt7Pqaf5ArDsHrE4Dlr
Mox1xuE9y7SwsUtZSRdNcOsQjQ77dLLJys5GvBseIxzOzteuJHMZJqPRF/DaGbduoiMGa/0KDfSF
y/4vEMqjyJ4HIt6QyWJD2MXlAHqQ+ri2dH3j/Y9PWywrsoJidBv/CVx98qkHdQMwlQtg1D6fUmkA
BS+u2d7BzhNdmK/Ozc4V7Xh59TTTEz0DuMp6x26bkcmv0koBq+E1Bg9X/9F69AP8J/tmjxF7IXlO
aqomdP2wHuiAxFAvKbqmdFxBb3FcCa4EkttGo6DslGVkmwf9AACMhFnumDDa867VNliJ4ewc5chw
4gTVbdkjqOaMdqk0VSLUw34k13Wb0g+gyu4rj7k2yAfAJ7iPlXS3aFw4yEHv5titzKnO4NKMKuO8
ucEFRimuYLjWGVDWQjJeMs/zkU6OJVacxDiKCCQdTo+4DpdJIAXxBezz1uzrHihCCBpfP6df/dY2
76mR1Nwp2FeR7W53jpNRzf6IR3biFbphx5KL/fhqDw5W8IohlRZRHPgb13IsEEkKlLndBWP3ZxPs
CEz4LVk0Tj1ioV8kMG3ADwDiQ889Z/1QvA9nho0xym60ZsIrqX/Z/YahT837g+xQ92u1XTVQDivZ
6vrxa4QDIHnUCFK70PXpPAAV0l/MFaBcWf+NXS/Xv6ey531/xSTOce16f4GFpFVHgybnkoePPWBl
KolanFExDXUD3B2xp4Omut3LulmjQ+83aQkI8+8zMCjminL9kev66kYOs79C9ZVHQ2o2Wt7TyoTI
LlC4ZM7Xchs7pQxRgfXDmOxWmYf4Vr9LqIYIcWdpqfCPHK+4fIYivoOKpzzVMlmIy7RnFE29yjbY
rmwRoezuacmHqhV1tx7yN0HLhhIq3mx7SekPuAaXM/YMHOSkLJ+MR6Fy7jGhpV9juUal8bIqIKuN
L9+L49MkDl3o4Kx6PZ/CcvaNN9EKaYkTNy/uxnIfmyAxYSX88Il0kt/hgJ+xm0/0RjlYMjyRr1M6
EhC6L+fVgTqRMSRUGZA9VmgI1IByIVmvASva6YFr2ok9wSMaarYGOOVwxdw9Iau0oVOIzugIXtes
RsP4/4gFFT/asssKJDHcDK3E0Net+wD9kpxBJG3qooiE1ExtMPPi3Sys5dfrCdA3Wqa/7HSF178k
k/WrmrJiusOGUQHjIZdrGFwGsbyuvWgmdTkojtu791eQPOvp6+0jBx519Zwk8JP3tWtRKZaHInZu
yIlvtbQsOhIzGbnzO4EqyWJDmNm0LJO0d6myVj4Rx+hv51nsyWEMULRSooWmR9w2NEFgMZT2hxqK
U5r06cTHNBlJxGrZEtxy9GvhMGti2FvOsa55ySbqYb0Ygve6aJqUseTyEcBNY0WgfHeY1EGTLB25
V9VBqlPd2iy65r9LWKgBKJhfjsoaAx7QhIXIOuBCXEn3BhCZ4th2ltr8EFpIGWJIVSAP2TWvCOj8
2p8RLmBK+aE2yCehT+tgkJOzCkSGnlPcJ2iz+BhCjEYfxVMyct7QJIsgLIDQF8+Wt3KdI2IbFmiL
5YY6vlbrFDhEwTtbfEVDS2qS4GJ1JEDvsRAGLr3e3Ixq6cD4GE0/1qPmUXOZLkfxnvpvhPEoRxZL
XMiHAUN8y9j97mciRSLdNsBvOq/SpIUwv89k/WmJNNBM8erdr9JY4GvehLAh3SoA0my3jw/KYALk
pwGkPwm2lfwZk0Nm9pmN7gfwK8uvVoKjdNQ/PjnU3srR8/iHTK1w5fVpUqv5R1ZP8zRcsnudk1Nm
p1j+LDxsXTRte6Yq+fGZcGGODwPypAP9ejUBGpYeixSuudaqmI691vYamKHCXOAZ24hWc+M/WFzp
hVEr44fQuDBGuMNI5XB+lRZPnfI7VDf8ZqL+oLUKVHZwna2f/pnzvSEIK7kmenREq/vAeZzmpI+j
jMCGVtXmSBjuH7r1a38HeN42wv403jhw2EqRJemyn/oKL6tzw0rHHRLnJrAYvUZYqrg8f0s930hH
a8Tn1/yHgFgd5z7AW7Sa5BeOXIyFAY54TR63EiIlg47/DPhoMc/pADnr6AKMxAvoS9G0RNupoXN/
y2dtGMQkRJc0H9hwjLYD3F7cBmrek8QD3zV4fZXaUSUT4KLMU42l1/SigOn9W6zmoL6LTlK+UOYW
B0LdaWerFCqIspRIIbbD60qV2reTkZ4O5pM/44T7C1CmzKZDtTbRo9VI76jyYESC7n9WEgxhfSGF
JGRkEipavZkRuhxE5WtpS9LuuHgz95SUty++gpOvFFLt6jr626hgqvqOLq3DfqE2O+Y87JK9QyYH
+theuWNc6Vg2Y89+uMQ7P/YJTORSLncyXzTUGKKgjNTkLyLVD6T/amP17ezdaUDgsk2YMLG7yqXc
P6F5BRkeSD/rNdW1YqNy8FQC7leBfd6Rp7v27XhseXYWul5++JNR1gTL/OGk8tXJa2M5jkuWmM21
i9hnRPSFyJ/MN9PCJxN+BjyMtWF71jJbYJ7iHbRHn3u3V6nNrDpJFIC2CBl78dob/UmrudyTFxw7
ANMefztUAlhSaMRiE70Vura6vl3y8GH57ycKqMsj9RaRISQXzpw5kw57SpDeDQP14sMmYhLlFu0+
DPChu9fekWHiJw3mzZZqiLUskZEC6OYRRJOycPkvFqnN0KcjQ1XYkf7JQ2Ru4N7RyYKx+Nw8yut2
huDxp7FtJEump3QAi49duwlaeFHIQPne4Lc4Kr6gZ7f28d68Lz77Dp1gApv+KfY3mZ/Loy+SGlHj
n3TmJcJjAx3JD8A2bicovDOjXsnB2Pv2L1H+p9ciyoAqFepVRiX1fWKGz5ge7bfxmEkrr49kUIrB
CxE1dvHx0c8FavmEOH93mbu/ocULHkmA9lpKIgUYn/PSUacHLVsgt3gmZJXklWdxsQB89UmGUBK3
KuTio2bL4687OPJS9AQCABnz0imCsL1JlkPMIMOT72Wul71KGG26A7ji/chhXgzcn/ZFFYabPETa
SucGfQp4/RzVwKk1hZmMecpBWWW05AhdhjUv8WY1M5zYXaRqIu9nsidF5LnaUxd3OaVOuPf1Xmff
95tDspgJcGEJdxbkQz0jrOyeK3Mms1fwr4M6mkV0cfI/omkYz/+3m6z07Reu7fc4+cBaPE0hXscL
AwuUdwjhs2mRJpRRVQvrOVg51jTEOQqNBrAOhlAd8MlFXyH1ZLqQFgOmTQXeXcE6/Rgy54v4FR4S
pDhulqkdbxGTKjIOctEk53tPzYmTlWtZxRDphcDDtw0TZqVOoCWWOhNGmXUjUnjVCj7dOIF74fQI
f8C9Y/M4Ml4OiuE/8B9HBzfJUS8JF8pviferhZN1vjsQRkVtTxqTPFgSYyZfLQTsIifAWzGwYhNX
z6w9qk2UI2cpToa9hMTU0H1t+EJQTt5NWyJrFQLaSAdyGgX99bBbapdtjTIbsUbjNxxAgQz9cvZ8
S67LqZIW6QFii4h5+t6257igKs1NkHgaIEEXIlUUlI/CUDk1qcgZJyUz2ooU9EObPzA4aFfdrjhO
bVrpNv7tFZuLgMrfb+NThs6ecUE8g7AdoqovLZcbLzAiQn5BloKIMP2NTptpwwy6KuAUbNEP+ZRJ
meN3sYne6NVYH3dOT/OQjYHYxalPnWADkpeSt4g4zfYFzyWqrr3hH0aNAt9CYuuj3qdlXQeAXTMx
rv/3q8MevmK6xZBqI3+QZJBK1GHF3krq9+elSdPnnAmcGkI4YUwWzD6ED9HMB1B61usqmuYVZDAP
uF4/o4C+Yowu6Fsyeaqwe73pDZrHMb2R8XukS91mofN+Fgudz6j+577XtgJe5fYycvNCLw138Kee
mq50la+GRXAjB34I9jRhCtos19rhGizRLY/LhJtlC2k8NNRtY5z4Ke491jtc5pS+uFSPeyMhcOnr
BQeAQiYLnaadFAI3PZ5vDWOFktoIJRgmUb3Nsr3rfDId4ZxYRl36jzeEUnYfwKLnizRaLRloA/9K
gCc4rkPMn4L4a5o4zaqW1ZS6LTeosYkQbsaT9VFkTMY5C5vXZm26WeeeGeRWdmmyvLjDz9LcKYV8
pDF+gv4g9/Wiv/zSXo7oA+1KWdtdvjd1IiBsXRM+ovPhyL7yoo05NftyDxIt/7UmCuRmNnyh5zoa
XsZcUI5ypJndPHLOOH6pRg1iBp1rsrTP8JvC1DglYYCAU6n3QGVMbvvn22mzJsNnR2KUe1+dYj4o
Q0oZRTTEfF5feJD4HuoStA0icHSJeGYePrbYqL3R1lSpfdnaN5Cvv7MnMqN9vbZkv89PTxq6G9+j
A1pPp6FDcUoHUzT6q0/VpU7QxLAZCpkecSbdbMNjMBu/5zD1HrSW9S0iABjD3/dXTbmjLeK+HR1r
Mcl9Pm/vLOoCwEP2R/SCzYnUU8B9tsEhoL8/El40gK8jG9d6ro83gHJPYZaXhp5kL/0ePLsptIqn
/YpuzRhqlyxq64Td0fORgRRldtvFZxbNgAauNPS3dutxIgZBAwQNUsjmB0ArsN0Ry//NvurNfkx0
CKu1Dh7NRiemmQ4FAptuKRhdoXTsJK4+1GjR5yjaoCSLmwpEE/HihB9kHR2WfJj9vBgf6anMaEMj
0opW0Op1rQxgTJovVp/culdoRkVzb+F2u1QLupu0JDXvC1R/NBp9iFkyYFzvfA8o9a32LwA6yE13
sv1YzQI8pmUsd4rzKKVQS+tefXXrB05Ni/a4RiG92rBZzLG7UXPaogbB5xynu7SyddxFKIVLsCDy
sKOH5nQaDzrBQFlRQtY9UfBbXgZJmBZkxBFCQxx4hjeUmESI6BFEHuPBG6jVQqYuvCZGwxrJt/Sm
ghwhQtD8tOU0D9lD0xDZ7hxjgqDtAMvswCL+tlaF658FjHTmeZSSIyTBDI+bhs4cOWh8BXObsYMW
J5OaAm1HY4zE5DOwhk26k8z3DECLC/5Vyc68Tsl6IoxaEwHYz60KuIfCKBpIe0IhYmjmpnSiS5QO
6apW1XrkSX45rWU4ScWNNE5Gor5LhI4+4ZXrczWkCpswz61xU/tEF3FlU2rDbir8dVBWJLbPzdyj
qya6l1qyYD9jLQUhEpmrYxnw2sr/VA7Y7AbNmKJK0yWUOKIg17DpVv+87Qqw4ySxS6bFM4buxWoD
L1mRGvrdZ9NNTeCrhLpiQ0Bc3vTtACmSRM3fZJZtV0TdhaaPS3b0pBAk4s2hUDfJ+e5JEoErFTV9
seYjZpmJSiAKwVse11vhZZ+yuOCUG/hnezJZuv6T+P8B1c01LRxehYQd/WRoepEyewz3pqY1TIEU
hF3H/Mv+nmPXhyNnCDXLNgVrk0/vspQ2e2aLo2G88mzpIQrNh3ykhV6Sh7KoeTcYWi3EUR/uOTSs
cB+lH1r76Of0SYn83SdFPzsm6sM6J8neOPErSjxblT08xZWusyucExHslDKnL7rn9s7cDsqURNIg
4tZqQv9T2I/8AerG2Hz1FpqJnuP4bLx9Mfyy0EcNWObPFBhe0ZwdpaBkmcI6qZKlxuGdN9MROKcr
7bgsFfnWyxe6Tu8m7ud2bGjbLIsiTFBVei8/cDwC5xVi6u39xAwY+cedqMYda9xE3omcfWuH1B+f
+Eztf0w9zN4QxLWhpT0GbmJuSRRWngTyTVDsB/HRQvu5vKHICHTjkPoMy+rZVIklYiQCDheDuG0k
o8XzJMP+gH1Bvpb7DaGKNpOjosKyIcj/uLLl0xLHPaRKy/B74vO21hazb1zrzghZNlzIAlCknNAS
sRPAG+dKDXZuz3hM7ObH9NxJMVM/eNs2iLQZcIID5u1dtlD0hS7JAsdcW7x3UVXhyaAHmYCqaXYt
lLXtLrC14ENjMeMfdiMN2JLLEJ0EeDCdbDjFZ+GYryVjKjzWVNNHzw+DKqfrv0SuEt7Vuwj09gnW
/M7O2tpENPRfrLAUzemzWbqx0kbSHMjC3ykJB6XROkZgw8CwQR6gtzdXu//u/jiRkPHLf/8KAJQP
TEIw36lP/szh97/eVnVXj7IStpga7Lx0Tq2ya15Kwn+0QIjFUz6cJmkDKaXSNSPZOEmUB7OGpaHw
CJjqgwNS5b+TLLPgL5IT/M2HZ045KOnE+tELAsUSSHMTF+ki4r3ka0sibVEgNRdcES0G4+JdHpJ2
2o0gtpYpyT7nY62su4s0JKqSAeAUMLg2A9YDy6ESab0h1dU/Iep2u/lNp7SFwF79BD5ErxLRQYn1
Thr+E74DxWDxRn/jw9G/VnRlas2MMAx68ng/VXgAvfSDDyyHODIrKomxa6woJdUIZ6VxufL9G4ur
bgq0D1r2ul0DadoCb4d+Aw4VqTCb2LKi6svR61/i2q7WkDwPoDIMr4L3eluGissIvDQoaSbMGB5h
eh7gfyL0qkT2svR0QQ/VJDVcnaUn6Jjeg9YVpw2PtZzHsw2frvh4ep/FHizhEMlYqcG8dPabPbcO
AJSPNJgINHBqVY1TVzRXBxP5N4VnXE24P+sw+olZBw8QPlVo2evjaDRCTQAayfMOZhnVNmsI6UHS
cY+JmSLZAwg9+9ZboW6gZ6yJUOC6fnALZexuWqKtHSZf12Raarg7drEjpUQGqGkByYs1bgzizpvs
CaS6wtbXbyGdTEAXHKHenSofNWgMiRSb2eX8nrmUvDzLHnDxf0yXnzLnqEqsFE/GcZrWuiuQ2tjV
3ZdU7dw7YmRYooEZiKfBg2Y+yJrGcWyXohHmChxWAwhk03kpGPB7pueKoeK8mYRMxeghmvpuJa6+
ovO26E7ex0pP48Zi+UUUZtM0LEzW/yIGEbnVunx8omXt6QFBKrlPGFd/EOsYhdatVqSEQDm9J2Qo
nXwznkD3z5AK70aScSlJXUdwFzwEXvAilVFGSTv0WUIbdQoIWdL4HShd4j9RZeGPGJ+GHscqqxI/
9yl6/PPcN2HYWzpCpUX4F7ZlUo/y3GRHiBWdqwRjyKHz8gwYqB+Qu4Wigh2AOO7nRM4/hFjoB/25
yhyAwD04S0Vs2PjsfvnnuGucyi9mMFaAR2o1qr9cUyYwic5lj6MkuFsj1hd+na0NCuLHTrt9K6RG
u9DTwpyx10P96ShyQ9nyqhuYD4xmMkjxL+/6G0Pxz860hVhYqJ8dq5V1k5nrD5JmrfLzem029fdj
4GxV2ktklXjLZL6FxuJUZ9cY5xTQ3njPUBA9bLZav8EqkpNiaFkLmkpifeayWuLj5DgNgb1lOcc5
gon6zQxpAgeqST68n8CMQFqn63rZNL7+2XMrXJ6i+jIKwD5H6sSFb716N4O30C3LJf4tOc1lJCmN
QAp3MdiJBwPwPkQdTOleRkXlJMGMKE10KtF9xSHe9ddLlc5n/9QBxwhtj83v7zTBxKDx17jaRdpr
RIEkLPzUlzH0Z05NhOTSVy9YlPLWtQv7KMqymk89e/ufJy5XNVPO95NbmXsemkRLeEt1ingtqz67
shAW9sItlxLYzT4A6wFsEQLKyxTNkQv+BaIjnMmehg2wXHRWGSz04HFoLREXqi5P8qcofIqHiOzQ
aS2syW3SMQnjPB9br1qkgq02zLTw7FKhs0IrMtbDH8LMErWqNNq23vqX6KhoZA71MSrGNgHw/Vo8
+PIQH8fi+sXR4e9GYkcyqoCVw28KdxrA9xjnCqFdQRJyUs+LPssGGyn/vMjtoq+dSvvxj5LuLy3z
nC80csFoKoWVtNBCZKlKa1EX5ovYavlsFc73PgKM8hxSGFL+WjrtzruGRsqxgfCgibQKnGiOYO64
1waTC/VR+R8zmcB9pajodOCvDnhHpkdOSFZjK+nOQHFQPCkOznF49YIIjO4DjyxULVBKr4IwywQU
2H4tkgft4wWovjNnn742ynktX2qAXgBLOoFHkrogwczWPjfeS1EaYZVY4P4gr13I2sOlu0CpSdPW
iNqArDZHsauJ6dIPe9YOhJ4g/8Ln4iMq1ubvFVRHSwq8DvdmR0ykodS1DiryFBfVUTKLdNPIG5RM
+one8HT0A/Xa08YYAMRsdJ6x+cqlEDMT3gLFelyAcHtUybhHgf/JpPcZVu5yWXsqRWLEabBuqu6u
HcJzsT9mPflnOH+sEYP5ebJ85cq+Na+edOyPF5dhwoZmPlM3SH61dVYMFWdwJFl4FUS0yJbk2u1k
sXUT1tQIeFoeqVNpVW64YzZbO0ryGQg6pggUP0JqLjTMmefYH3CSGcqUvXfFlqsVA8hHfrbPPJR8
N+ffeGQk9XlKPSfVu364DNA5HD2WWaNe9I4b8cJUxtBS3T1ZqZoDh7hfqWvOdnHK/9vJGZP3V1zd
BVfXy79/K9rESYiv+sheVcJcxnt+JUuz0aqHhVqcFAu6qM44Q4eGbUPS9ocsDlNgn5Hv1jTi6sN5
O4svl1XC7ZzN7g5vOXZqG3pXgUfxxR+j/rmX5hLTl3VdcAHVD17qGNzTzIAPjf8r6RNVs7i+HWpO
Me7nL6iJ8vlHqi4JyJIkGh2/0yVFuS7q9PYN91HIhkFKPAVt25Ctj7xFCmzZCsm3C2+LqsYXBfWb
sFUFoRp21JINbAW/mU1VFvbSoPM3BDBll57jWFJw/8ElIyREDNeNWdumMRnaFfOXFAKHts66gY+m
l6k8mKZVbtl87PH4Ny8MNeUGtYCi+71Gb6mxdf2ub1ckW/oC3EHH3bc1BRbE1cIfB4VWKtwQPmkD
UYXORoR6XIJz8aKqLT+4Jv9UYw7p6nEr7QfIpIcNuRNYAloKw0LFjNfW2GK9yX37gWmH5nINeJUA
bh/nR+qc1bDTdAC8bNnNuvT9phtPmMNMM92TjV6VF9N3AzYbzz8lqnZiFpBIy5xfa0uIc718dtyY
yh9PvEIz/lQl7zxy9naAXpjfyY0Uf4JmHD05mdrh99WYnA8nNMiX6WuL8p2PdHuRa9iLODOym2i0
iUwCALdHjceHx0ADB48fW0xKjppkwHH9FKeU1Vp6/jKd7XfnVZSjyLMGnmgy/ohngV8zDQ8erWY3
MKAIg9xI3FlPBl1xFOYQYar+AS23O3ZvqKDJ0vcHr3LevrQQy992LuwX5zIS2j+PuKAJLbY2b+NX
HVNfBbKiL9Dz7lYczP6i7C7OeRKvfQRjMcKfgTdj0u5/H2VIZOIwnIF8sVGpp/F39W6nwPVj5paG
rsOxtZGlp0WE6pTLNEMjwhmbTn60uPtLMwkt/JVQMo9uTq/Tlr1q964PSTAvctMVqQ64aAsxg6zs
Bj/TxlsmxI6uCpvlWthSgkD7zB3nt7nU/JLuKTJlEl/WvCykQZcU1h8q8xQIRxwczaMGGXr4jRKx
iMTFsuHZmWEgKn1uQCTG2bPAh9+EghpSbrotD0FQcJPl1+IPkgvzna4O7RlZ/j268IB67hnUI2XG
hux+jD6uo+Uadze8XHWeDHsW/nABL6IyWDBo98QVm3FewX5ONL5M9uFMcSElUSY/Uonz/xZ25scv
3JmUIDtUvEM68rFVEqqHDsYhx/xe32CqLy5BVwuwiKkwMzmVEaB1FnjK1jIKEv2xtNt11gGkhamh
34Ue5MUiJ3jV6ha0xbGziz2djr68CxWh4r0i63LmaSN0cjZUZl/5tTABrIO3Jb+uLEIIRF3sA6E6
p8KRXcYgUavM8/0VLL7s88SCGhJ7ANEZxIBEwCr46G2N0YwUPN0lu8uiK6G4EqlOHzN6U3ukkV/N
HkLBLndYxENt7DZ+RfWOyaDK2P9kpsVsLOTNzdc43LeMZwVMHYjlN3WpNRgahdi/4ipdEX1SmQOG
Ww1ASuV5aI5IOYkdH6SO+Z+5YpEyWM5mA+MAs4pHt04kI1/eGbAzpu4SXwPZG6O4yfXUphMEg4P7
1xvZebI49Xmn97uONtVSWogWNywD+rJOdOLKL52gHUaOh34C+BXbpQj5j/LTv/20jQLRU1ZGznHJ
2+5b8qowjEQU25aMDeZeeetedf496q/5l9RigcyEr0m2H3lCoJZizAiq9UkOOmgEpK9l3tR+7aj/
UVeSCT82qb4GM7wDi1W7GuUfmfGe92r1DiMlc7K5RYRec+xCOqpFrohFeF3Fyg13hXTfQtMKTU6w
21h5ip7aJONf5O9wi9/YJgd1IiX3713b+bFBxyNriSJvhJYB6yKjLXKJR3J331gix7nUtfCDrMAS
EK3PfpXHdVvuHla8r4FV613ilqbUJUUroocTQ1V9wmQpYyPGyX6UN/7z1Lx/t8x9l/Z0F+TksXxO
4QgRoFBWxsBf9aCnJHxpn4KvEIHWFs0GXOzQ0DfeaO0vhPt50u/jgvQg5zW7By/MLBYA0TOdVb14
HcWU5Yb5GfPuUuA6chckzsrLBa5iwbQm3+s1qxJeJzwnrStKzYAYMx/tRdafMVDJbvkMEJJ6G/Tr
fRJjnGbMaTOVRqMggZfR4YQruEHNUSb9mdUafHq0sWCK2cChqTLFzzKjGVoXEHqeRR839cTW6PY9
NZcdAI6viZWOMD9m8esiDN82xenSf4CBtkEQHdXeqUNEDbTdel36+PxYR8mcot0RvwAvwNXpZp41
86fc4PXoEQBrU43aL8QmK63XLC4QDUreHwGa9Yek1vuzGRo0yM1SnJWtd+oJoxAGguAhsbNxwQOc
cy3dCyttq5GW5gJSMKC7VrWd5Mv9v07U4KPMcF6VnNV5bHZQv8tCHs/1Oc/tDMS2hvfSNIXg7MYs
g/XC6y5dZnHUCnx62fHjLNH/wOWpt52hZYj0dIN5GBwciMBEjLvBYoLJyJId5eQhnvAn3AuhTPSk
8mJR1ydq0MrUowcnrDTkKpv/csfcT087jpmU6bfFDQs9sCxeCiv5pDFV6zuvLAfx6tfsCRmpPNXF
6yZp5BibyEHjkZfaQE/qPltaKkoqpvtLFsfMZsiQKRfDuUra+yD+9/xESGYZ59AhxCIltsoxv5sP
b5N7S2y0HcuTt/jZIJREPFYbzj3kgYBinsAU9VNlkPoiob0VPKRyIjGKTvAck+bbZ1cfCfE8ksCn
0eoUEtYcLONSyCGv/bcG+nFoGgBR46sZT35+WY7VHkL3/qwgqsNpbA2Pd5j995r+f2UAJB40XAOl
FGN4KI3VnZFHL7hfEg8TN80oLYbvH/vK1A9UpfLPwZXxtPYLwJDGKQu8pMOhmefm9Po7zc6kceuH
3JqyE8pjqafaZbACkHtEnXnM3ZhOnuFdP/JpwSj8OrsQX6sN3Exa/V0w+ZlSRb44qAr6jKe0CAhR
hC9rR4bf+kmAxWrzAmqgNXZ/TkBEMXghC2A7AfWA7T7msESynctzzVnshchTrKoXBG8HpiQyDHY1
AFwc9CvZT2RtTBK8bhtVgoKeEjLIRmeK41KTqAukPYUwAauWdT9Ujq1/JgSdm5u7jN2wxhBJoFdz
457UmFoPXh58FJv/8eqEzdwuQS+12ITal8MJMQSTyhECWn8x3j0RF99iFSTZ72t7QM63JCrImAUv
U9EL6lhFaAiY4FTzFbsgbejVjJG6Zc/WdtBSScg64DjF+mFRUegbVrruQpsAkxfSW+1sYGnwtygy
boPlMxhgW7zyGzg8T1z7Wrr3SOBBPa9by7pjE5CywlPsBA8JMNQlRi7xb8qEL9tNZWZG5/d40+7U
L5Reb5T71eceM/FONF+KRsW/3g900XUksHXOehgsBMhhXYQ4TxfT+lW7saEdPL1AYFqxXjmIHh9g
YJutCK5IX3xSVabqFUBuZ5BE5jxZSPZjxw86QNc+ZBdvx3ueM2tNTWP3lKT2NdYJBYNlJrMW8Xp0
g1AiwdVvO1ZkcGKnOxy7Udi5yk0N7Bd0a/Brf66bIV8gx64jDwqaAc0SdB3SlsjlGQsbTZGURy4Y
XjiPB7/nbIR992a5qbUsRc6VcJ3njBJZHFwP7OBqySSoYJO9YzyTLvF6KuslylY6asDn/LWHpp1d
ntqAX1YHPDnDJ4V9R5d0Rf69q+XG+sohzE2vxPhuCTrB7rNu/j/84HRNPcRkWCPah3NA1+pUyRiH
A/3Z8PgdTDXnp1fJRQFnaykz2ZmIgttRuN1EHTLapErP6JfTFNZ+TY/wmnyTaciKLEn8q2AbBCRZ
0TuhAbs26KMT0/6oEAo6kpzS4c28NwuAtS8UfFq/1fYuAjoeuO84YHcp1ito2bJCJAesFDh5EgWg
DQY0fyO+HzG5LcGjJfpNeLOdryfUheRagHM2AJgt+EKgNHIkzlQ5Vx7t6NODhZ1Kv1nGWW1OL8/e
7PHHp+86RxRD9j5DF5mXREAAsM0hYHu4j9oYSUT0VAPn0K1oh9dahhieiW6sJZOfmxGQL99zp2GY
R5UM7/W7vq1r9KusN4RvudJb999hwt/qHk1q+CxaLsNvHRMcbhZebjr9fkyvzK57AYxBfrMJXkts
DPsftiUg6Ff7I7d5FT12SgqUT66rJF+G0Ny6I6T+CtKD5VFtIVgdyr9ICoGvwuo2DWLxmZ6ta3kX
KrbvIypFeHtUp4rdP3vbdnteqpuqsYl6qye58m6kPFZesc7+bMigFFisN/z2HoAUKt7R8CmGR7oc
Y+ZUltbQvdCmRGoMGuBXebSJbWOF8rfy/UCe4zOCFQTNeybSbf3C8b1U1dYZSEc3vf5Kv9vtlxGl
a9J6RYkdLEAeq1CBqcEA6KhFGcY5anmH5hzqIMUJSnDrbPIzPrxTaj6NfQ55GoWExtz9nuTjkwo7
i9iFc+cRVwl9yCLTj8CN7b5KqqXW4Bd2+rVwyIcqUfHlkPCHYxkOla0YJ3ZTCnKeqlF/hHpyyhld
MHhgGdTiNlprkDt3tlZYhiEJRq0HGkTl22/Yl0jpYBpRPx8W26CikBK6/NPTNRo8zETcDT25pmGC
amavQ5ciWb3ZI9QXsRctu0bu9GdXz32qm1V8wINjxO2zHUZDr341TM81Fxddmfu+16VwBtI9jG7x
1TE7lqKUaME+uErQ4IPUHrWFcN4xg+wa6oc3pasYUNbFvwDDZN8aUlvXArPPj93k9qsXQ8Z+JEHW
G6tEHU3r7QU+Fo1wvDcT1+aQ7OiwdvRpwnzhlZ0VZndEi5v8A5Dg/XDc4QiKfXjoLZuKQ28wKS7L
whXHnikJQ5GAW8sBLwls6MC+t8iENpc+GCFZg0GM3vjIMroC/7d2D6e6UOv2IGXd8JhvKaC7DTpM
c7UZigehI5uUkt3LgSkZ54pvw0pFycG7R13GXdT2QKxTLoDYSRizJKBexcx6Y3SauhkEvdnA+ypn
uMnhYPugXwkJBp3SaOWIR3Z6aamvI8umihF+RIlPZRhiCWLDlGp6zGeBbLUNjEoXxkNQ7kTrqWIH
iBQ4n0HvjJQTFCS7kxpt0V7hilszc+Rhdz6orsAR8PkRT2WfUy9+hRRBvP5MjNvrFLV8j4mZdrQs
UTrOAsV9CVnXPsfNmTAxfdyol+QnD2ix72YEU8yzUdt3zFs8eHfLu4ITdgexyZ5ayHHksU9XaTCq
Eq2y034VXNp6XWn5SX+sAiTZkCvJmLYsf1fl0BfT7TqXRWm/459UdqUHyIGQDU7+IPZ+xrxqoWQf
M3ximSXwD3meQDJndYcy8Ku/m3qOiYseuCrrhjFebjEUhL4Qx3saF/KAgPhE0+HSIEEckgHM4Zye
vfZribYEGATqUvCmku/KcWAxeGLFV8KHkN5UeDMvFfSKr4v9M+SjP7305TNJC5A75Kh8jvHyDp6u
u5AWioclvv0UzvjGQp4NNPWUPe/ML8VeX/V3llCQT/a6g/b+CwJUhMgXd1c8Im0H4ov0rZOQTz0N
dXnuY0nC7cLGQo72tffIelO0vXSThbZYS2h/JdrYfHselgYm+K1T3KtTtkGneTEENmwevOKHzJRs
CC2kjvuwKNtvAvjOlNo9K7fphLiPx7bJTatGLV8Ebx+U0Y7HaN0uGWj7YT1AE+ICsuR7+82Rg+3D
Dlv96BSAF2HIi6xbOmuSGslThogyfLxrw7rcMx6O0Xa1ffeQQMFtRV639X5akfvJUUfeULaHc4NW
L3iXhZUvZIdRBQPM8UpuxipUB6FA5mYE3RXglq0zDQAR5u90ODZBJ1kNhmoedXSX4X84tE/P5Gr8
IVdNufiC1ewUpPSPRbv0CAu9+bBAfAouC7kVG6mHyv3QNLcTaFCawTQO9Eofj8xXc4caiwPM+/3Z
zsKrGgnyKXMh1kq7a5KLo/shh9vkcPlxYwUwbd4EC5izBRytwXiHr7MGOKwcwPM4VaVdo93U2FRm
QAPlkwa0KUmNYdsh6DBjoXFqARHS7SkSR1w8Ni1gxT4rp5f/BEMvPrjFAdcPdrMsQLag/+dvsJlW
N1gwzxK1RcOyfBbu1ry+F3Q+6Q76xSwhe0uGu5vGCQ/jVL81XyOjILSDil9SYoHrgVHuFvH0BoVn
hjhfDE5oMNRBR+m3oI/Rl91dwQFupyAHAfO5kUQ4EQkfFcTAwaIJiK9we1BkSSe8rkmHMu4fAGTH
W2aNvOrEmiCC1Fnrqhe2FbRlb/NgOzSVwu1yMdZ0VBHSQD65Zktjs/lVXBtSAztkc54VIb2GCAoR
ZL4DXfuVSUqOH4XBFbWUb+zrOaNpUigKKrk+GxZ+WK3ioxt7n6QFYkNPlaoSQf04I6bBq88t7KBo
eLVbu7GsRjI3WAgYPXZtDfwMg4cvhwqI+XIyDsIDeTKV519tZltvUTINhSfdy5dORH30wGJ87dP4
i5GFcgsPV7YM/QV2l4Gkh6IZyesBC9ScjlcHqMEnj5TVmiSh+LOnFA2KEW1K1VA9X9KZpGbN+91s
Pc/noV4/kmc1/HNZmFghbJkmFyi3dC3OGCRNxCtDxr31wBOg4024pcLwF+52Mjxc78uLyw/bAfGt
d0UzHibbfQuPshAj524k6sqkjFKX1rW2HKTKlIYK0878F73YRs3+lM2v4l+Uu+bpKc4DytSGwKJq
5BT3t8Gh4a9MCyx61UlSYQGCltsnq6g4dQMMsZVcNtJhzuj7jDISsexb8HF5kup1hW2jSaSuXkMU
uYM88Mvz5Vsah95AQGp26PRmOnEqFFICNPUurMTqt+A+JcbmapyNCRReqXj1Y/NE3fi97nF2LkeI
k7rcS7gXEu36ZTeT0qMLIlbIgZZ4zhZIUwwIcabG98hXMfFSqq9qh+4xDngEp2VIYz659dI2vNd0
HaUsete4WwQ8llPt6bCdkCrN0Skd5sASgaRra41Ee/eXMED8bhuuyyPajKmrW48muhLUHUwB95m9
pMuM8z5V3Ygk4iCsY8YRNUtFsqtM9S8G5bi5ncthG7XlZdK2xXwZARY9zSLS4ZqgetuZoY0MC88/
/z9UcP5FUfypwuls0kTd/zMjTRuC5m8/hhy/+SD/3geiN07NLesDQD6Q64/Z17vvvOscM5VFV8Re
DUQpAjAO0TQKPbkiyqQYF53XI6Eiubkn+QP3NQsGEbIX8zgYTCXYaTq2/Zyo1GaOtxhlmAEgfmWy
6xcv9uZbRElhTQAVv5xW1yX0FomG6VESm7JGWyeABW4BRjGLb2rsMVNUI5SpFggVobRXFFSVRjQ7
o5bVvU8PpGuHtBZKlDwU0YtG3kT3DUdxPA57l5mMzECP5ndgMVMSFOHg98MNGyi5DJmbTPdEBwGH
PiCd0O4tqZO0bjdL3sa46AMK9Ew4cJLF9pJjaU140a/7eT5XSNEZSD0agmh8KFN7sydBDKJMLdNc
TfrwBqSehAnjGZ3T54cPBecbsiJaCzATL1fO/7gNl7fDDEaKndrYs2V0D9NasK/c48BsADJRG0Cs
2qPAwOOYQSs3oLCyXBjxhp5Ubg9kuJ6MHz7ihA7BOC6y9/vZlS5tuPnqulNFj+jUj0vKMhLaS3hi
jS17os4FiQG0H8L40okMjM9/dUpqdyY4E1WHkOsC74d1wRmzBoSJSD1Nl3wDaeKWfz42KZRuReOb
4YvSI6huP1uvp7FU6YZBjspPdLSryqx7fe6r87zd1x55gOmS2AoEt9qMxPDjWq+VZdurnQa8Wb4a
xO6SvHvGFwmPxUQBH1rDOe+eptPQsJL7th4SKUDn0jhNL69GcxoPnCsFk+eag4e7HZrLxC74F0O7
hFjqClMdCudIkoDO1pvVHYAffwpaBM1geq1Bd/rjbOff0oc5r9VxjYmOCXG3+qfMdS2s20EHo69G
agD1dZvAiVcJIWFqeQtGrXd3I15rzSkle+trSEKe+4pKVtHykoIsIBZYdGtsftxw9hb6095kbYKw
U8ugnXO1clEvfqvreA3FyA2crLiRRW3br4ti3dn7ojSbJnGu10D++Y1efAqMMx9qElShBQpMhPtp
kknPtRH5hYgwkAIaQ3wE/wJoFW/H0mI0gXXqe7P1h8hTAIodBDB5wtfcomfOD6NYtD+I00KF9SoV
QnZsl4UPFnYESd7WYo/BY87hPtMivexHDFqMB7O6IREVfEN6gf64bQnYyH/hEdaVicrJzEnyzPCS
xlhsAjc7hc64sR3I6LvlRHB+hpyw506nSwOU948RMpDPp6QaRTXHScoaRIKoJvR4xVqejUgqs9hx
02y4JPTYtKV6KO8wLRQT3su6krHaGDte9s3YQwX55F5ooL9EuJhGJqs7G4fh0MQB+MkSAyd7GicM
S6iYaV4eab5VCMW/Kgp+VpDrlDc2UORI/B48kXmGNL5U4juFB0mrM/kKSt07iGrNAemY7/CDlqY0
gAETGyPwPQxehe8RjBzJ+zgEj9YxSxb85QUnKy0iEtTk6wKLzUL42Anm+LGx7qDZPdlIka6JiUdK
0cFld4JNN0SGRCS9JeWnfmjs7HDeUDA5IMWhbTDNsI9cWv3Pz4Sec4Cis/iI6esJw5nj37+6yPD9
mkJqgDuaJRNb1Yxxy/zwVU27oAxhVBl2LtDfgUWHEeU2qO+OVS9k+t7OIQYg8NbrrnjyIAjK9Adb
HwZawXU4pIUb9Qamas9C4dwMIm+8jb8dbWw7hSrHiFDkXxQj4QF6egyi935EoDsEREj2P3bUKbRK
G1zJoJg3NTo3VJkaO5iR0NXO4boYbWTON6hp4OENyp9983Z1VuGTxA9fEacChZZxspkjPLbKTw3C
yrIIE9KqC3FERhnXNP2sOUwznAT4xKXYFLLvdYXZadSRc35TEaKTJ3oOVuPFGMj1KqX0nWNkBZfS
EHTNUH4MidbgvK0ESc1JYdAVzZx6irotB6AZVbbHmTvYM+xBRkitLFsatdG1yU3EKBZKjxUAs+RV
gY6XXYtn+GH3rxbLxlqrY/se2aUItFYEWDFDCxkrFhGcp+rPrtcb9szgX3A5ZjcPZ4CmaiVGx1S/
Hfra6wi+Y6N0LjJ0iMXyiGb+HBOsLVxJPvaGHGXRCN8sDEXybz+S3VfQEtilQ7yBL+8mYQ58AAWH
wOirsSqC0xhmbTyDjlqUcnBv8ule7X1CKH7zBMoD2PVKou5lqAIUWbTYqttgfwjnfMCRZggn+2BT
3djXiH6k41Z9xy68/MTUgvpygre8I0bAJyKdjAm1ZZawhGRXOMP+sBOtWK/3lNH0d7pddT9S/e3g
a8I4L/6AU1fw5f9fz0kAracacqISQG+r53qOgy5nmeaQ6zQObPZVTDGUiujy+qwU886xGFpLNy4X
RtZjFdwZvVh1Q0r+5L9CRPWh1CwPFG5gT1PxBhDsTvPQfw/sTov3fTbS48SFwbWwt3nbVTw/QSm1
3qkDCVrJ9jlmCxYRqwDfoVtrfvSkTJR1GhvDOUyDfTo2grzJO4H0t507OtGNeiIe2TbGHbIxoU1j
fV84UCD547QnnqwadwLePRJXUbzaAc0u/jMjahX4z2Yi4SbMvFjtR8+9NPRpLp7cjPHugRchoeaT
WZYpNFVMICrirNIg8NMvGoSbxi5z2aakXTdODrb058b6lel4wlE68xAD141fgNXbVuVeJR7kVEDs
RKWFXsTtdfPnsSeaEqLh/A82ZgSArk4hf1PW1abGcWHmkfyXsq5+rER5QBK9NKy5YNSyNMpna8/1
Swt1Vk+ThNamNiw5FnP7ocmf875QebZ+lWGRcwkXXSP9aolNoN9QNmmB7oxLkGidA/gjU7t+73F3
N8n/0/TCcnQvHTL+KNliNYFmEycnB3QVmH79ji8Ru52uPWXLpyTkZ2DdFaSkMNDp7Hdw9FMyY2zV
IidMEVTz+c3Ndkr0YwsXF7JgOPEkMJczTQ9DAPyTDvqSHGKoo/m+0rXT/kCEeUMYUP2KRHD6NXEN
lc2NpvHPyzQXwnkyjJUPfpO8eYFm/IWdwRXkHaan65Z6LAccvK+kw/YY0SRRyFhDsiKvfVGWaBtX
ADHZB0XSgCSnjGInONB/JYj2F1KCfGgZET788gE4J2XQaysiTiwmuqt9n63VfMHgEBZgtzfg0ynU
Nb22dxrjNca8HtHwHUcMs2DUwZVvmtG3QfDiwIKqVGSm6CeRXDdl9FHy0Cj6P9cFT5moWS2/d1ci
FMT8NOtVmhux2AdUz5dDlxOHliqPxHE42p5iaU2/Aah6cMiJ3OWatHPGjiYoT75X+rpUuWzWuJ2k
qs4MVOSdz7mwwvD+KHFYRwE/y27K0ocong7Uk4pnq3yR89kiMM2tF5vbOl9klImJVb4e85tyEv6G
bnKgFMUEj4RyPlMj68xA2fqMbHBfHKLMVOx+OYhpR1L548fY8UogzeGnVU9EWwNAh48m0Jg5cwj4
T1Dw/PwTOwWlHuvTLoQ05lYmhlD10hJaQ3uCiiFgCQMqH1BkCMkbLKpUhK9Dr09I02CnplWTYi2t
3Cz0Jop2vSKmj9SCRSAjrUWG/786DLhU2r6Yv6yY9CXDzuLGyGDNlhD5iWBda5s7gV/kObHYA+Qs
5hZW3/pvIyX6EgwA93/d3jMGudOzoQg4IO80cqMWN5mOVsg1mSSceVvPXtYcqOyTsK1M13PuMLQl
ghJmhh80bKk7UqvRofNWqut8aieOBIpzLhDklZnjWjQmswrJqV+0DgHT4BAGksGdzJwj3muMQtfE
VTJ0F+CinYub3oScifSNvysOs+oHf/pYir0sPsF08qJG306q7kCa+ZgBMuwArAV1a3ogXVr8W2Z/
ZPSHRZYk5NHx12Ol8p/jCZ6sez2guXMxuNlgdEN8CIrJSXWSyCT0oM0OyL6/aOVO5agQE18y1gWW
GEogfztXgGAoh+kihU5HL1yUrE2Is7E2lNI6RsFthjbstEg81nrIv7KOVWDsm/Dx3uGmyZzoLT02
oK71GfC38Z3DnjLpx1tbV+/YdsnqvGGgpQcS1EVWTgpydZ7jfJ6g/kwgnv78Rn1Oi9jyEIcDJiwJ
cE7zu+DOuR1a9hBo/n+VxuTvKaXr+GjPM6Cu+hmro94pjE1wiH8BZ5/+GDZr6AGLq4l4dRjTHxbD
iX2qIuVNo74KTshtUUBFVBHdP6iIuI5iUcFLfZpTi/qhXdixVsRpuzSIxkViJNHeZJ4UO5M+DXZ9
mfzYISRDzKytG8fvQ3Ra7R+Cx1XE+J1/RUqMs/byAxlHgoOCXYwfxmBPeROB0xjRJIh+2DTJGOVh
PSormbvXxKsCVafA7020pJ7KbVhwup/iEjvcM6p7AKINprjI1CtJnV/yP+/Dd28Qd1kBiyEuJ3Rt
sGkLMA7LmrmWYBAPJJcMMMBaUM646hexyKn8nn8qJbyJRYtFyFv3iJUXX3a8ntDI0GHpzx1zt41u
wgG0as7y1wRCr9EspbBIWJMx3WFBSSx+5w0RHQ6JYTCzVzEbqMwYnDAKkXRp/OJiDPW+XnUZM0q+
5SlbQxyya7aHaYwkU4rYdrquP9N60mu28JDCCryS7RJG98Qyknsdr3OK05DHbv3TkuJVenpqyC2v
9LfbkkBkV0qVQB9BfJCukr+mrrPmCYJrW2hPPOebR/PL9R93kf9rnn7H3rgHiVzzVbltuaoLnAf9
1AG3K4griX+jPODnKfIlrAlQBhI0KyqbfGGa9f8iZ5Td3avOHO2b7+RdSrJacxJgJB4cO6xguUOA
B7PzUABhmMOIEWslVO2DI9dsoLr6kdJ4uSxGQe3Pe3mtMpnRb2kV3ORpG6ljXwIjF7WNSoW5KWEy
JF/HvZEjAlsb+qyFyN+fHuiSALnocvS2oxy6Y239fjVERH+bTMCIml0yK/mLIQWUA21dId1aRcjG
RdsMI8qrT55gNbFhuybo0T3BqpBRUt/rjNe/kfY/mnUjDvh4T0ManleBHRimFwE7y+abfVG/dJZ2
9hWDzlpt0jnkkYk+8g7/wzWlJeQAhC6ZH9mUpA2L0nEljMWfG82sWBDV6o5yVTUu6QXAaosOmRXN
4tV+Fik0PfE2/t1EHzBuh+JlpoYuTdfdP82/18vmo7iqoPROuD3uYjhxnibGp8yMB54cYYDPVjVc
Q43spgO7a+vYV193uEXhqlawkpFZfxcBMy6lP3RJ65C3j0MVZTXJD5Va2Wpe1JmmV/D/adyduv9m
2/Tn8KgpvGojNxO3MqaYKfs8nFOKVV6VANHLZqWGqyVeiSaqIAqwFivOyIE4tBa6xMdQx9swwM75
6jXQx1TszgU27iIDD6CPgAOIZYAz22RlgFn1D8RAOtwOJMI5KucCa+J5wpmjWCmVFfPbAwpY/V0v
X1Wn9B5R9XZEY8nFd6afaUVfDBbiM+L4eAV0/kY4FzBVc56P0uyoOnuUYHMNGoXLJsCuDTLMGO4h
M3310aBc1TEEegsuzTkglozl/guUDYGT/djcBURrSabPWufXH8C6IZIgbqyeC94mg4i2uZ80zPEQ
aR2SkVileX6t5NcvyJ7CjOkpiTCeKJc3elVfGys9ew/Blgbj+ECS02W+0iW5YK+jpEMA8Y21ag3h
azrfee94LcNBGTeJ+Mpf/p6R4dWNOlb4Hguujpsa7QxPn8n+R4TNfbbjdbn5v1wSevYVFrsT0hEK
O6iUEUSXMp+2mKT9uK5LOF7cGulAwMacI8ylCIn41vL1T0p18UdwjIBu9uLPV+CXdjFMBDV+Z/0K
JxKF2wDEBcHTIEqxRZg/s4dYWAesiFkiOfksWMIu9brDFnBCdzZuUJUsEPKWjBkjwVJcq7lSmbtJ
WAZ+zp1p09vS5Suco9ukPUe7kw91zSgbZgwLV8vqnkFcGk43MvYFpWh/gcd2jW6Yzt8F/9YrSCKr
y1vs6Oh4teRkIrqcTUG7qBfEyE9gAFOhtjRLxhnMGvczXNNqQtGhs/JgpmtvfaZaOjBnJYkBI6DA
oCqSi9gfmyIjz/4n6PHgUerdnV4wWehuqo3SuhmJRmkeal/NW3rjXZCnA3elhMiBcV6F9Wgzqk/R
Pvu6NBXeRS7RWnEDc1nHNKZoeX7ljSb3rpgIktd+kqRtqa+LsLVjkECUFOZpHRjyDrUc1NOQkg9w
ts/LicnCzg+8Tr+kzgbQLbnFTExm6twr+d+3eYiNCid2XJD4dQU8UrZia7wrOCvt/FYmzUBvMNRn
R+psJVnlAiSSdB4Rq29RiKy1fJgDE0tmAnX7qwlDgk5ViCObR9B9KWvbAIV5ni1AN2VACM+i2/CS
F9YHgdMogW19dtAKx9HtZ5hKXRpiIzOIpSdlZftjO82KqJyFr/FEer1QTCVINR+WEFn4GpM5RUY0
OFVeJ4f7iiZwj0tuNB6DJ/0Z0tM9XOrU2g2ZrAI7OIl1hp2VzFVUWrMERNmFZKWmnShQ3UEPsusN
4cpRMr2R7vKd4RZ67eDkCBAXMl0RJTEt7n3jkxsBFT8BAgNpNi6ou7vlExf4OPncAOtl7Tf+xdUv
OwgCgqFoNe+L6SnWaI3V1CzE5WcWteTE/1qT9dmtA86uMmMNsA7WgxGJmAjbmF73i4LYGVx6UKye
MqPELATttq9yn2sIqh4Fw1meBmdiSwzO5JmPzps7kvwAU4lw1BYia/krE9wMTWhuZD+q7q3+ovaW
SxR1hPj9pzG6/6dYrkSIpO3g+cO64M+W99vhDvobwAb86u890ylS3047wBuaIcZjizlea5GKvrBX
doxOb9YT/wS7MAzHbW5vZ2GnPI3SE4dAkmzWsXNFMzOfPPaMXuUKxp/g9gFjPKhoAm5M3RpvOYI5
A/zunctylW8mKEO8NsA/lB4ukQufI+iQLcN6NP7YqfEELbRD+dK2a4FVJs7W1qe3r3Cgsr+lVwjf
f/F1ScPT9kn4HIGAKzdJ4CocCTlsNbvi5GCoUeKzo5jsFv9Ix/v3nse6zFAgjxu/OprnQPyJJGyi
DAurupL+eHszf2SRJZMrzS1jWx3ZYxS7kcmQYclkAIET7jMTCRqYv8duFS/jt3VoxRed0winlzfW
CRk63ApKRwN/BQKjUAyKpxspQff/mdaBn+Iw6x/PsPKpdcsG+yrfrOz55ZJ5ejEKaRxBttyo1ytx
o/FJWnfk8DyQ1bpG0wq00qGxDmeeAoHS/L78guR8tOagoIYOz7slz2Efpm5Fcodvh2N4BxjCzJdt
ORQDJVQ7y+eq36k/QMJSo14zn9dr0rjN9F++7D0aXPnWwZZxv2uXNp+4HuywD6J9Vuus7lZpkKFK
oqq+u7sitD93yQtM51mDjanLHKyrQHiS6l8mkiWjBWQ8Y6DoWYImlm7d9t04EKTasvbdgP7V+5Ir
ghIHUTOMS+NPKByOYFW1275Johx6PbInqiEg8FtuWpgUmsR/T5MUjBIUShCDjO86mYCq1guU7lCC
uPPIy7TPE1OTEgnvDNKswttN3zQ/GzxBit4LYyQUri4v275lGBqa3x5czoaeIXzWfDQpodnlkilb
2hDAx+a8dn0p01sivZR2FE9UfCzyak+WJ0rc24J1G1LOrp4lNdb4vVZxRqVIQ/vSrIB1w7Zc6jus
x3D1wN12fJVp0nRVu5HajooRq2QWvtTClqAadNMtUuuJE48U1vExaeMFlefxA7a2Uh1pNYosVANa
5K1R9K2HUIptbFxv44OIysBPFAKh80bVYFmzVt/XZNnOrTDyWwscnEZIvKQodX3rw+MlNz+QjgC3
azkXNH4ICsO9FgeHb2ZJ6c588hPVU7xRQDvnXs0gi3+aOkkGbCi1gDn3+aD2NC/WqLoomoNmeSWZ
E58zewv5LEjLR5sFseuvErY8xhO9DmAGeO5usB90iRs8TqPjBvl4m0FRRr/9YuIRcnc6rd+Jnw8K
RoA2oDFkIVn67itbyhFcCi19nCaSuckGtV7idNsAG47jXvklet/E/Y01bpgAjFYKn0FDMeJo0ysk
siztxQWcD1BUonsepOYIpZGels4AsrWlP2voJSwzK5Fu6WaZkyy4ohcF7Wzk0BGHg6Js1AXoIQnJ
fiXTMnL27baM1CdbHcfCgp4IgN+NxKbYanjyTjlrIZ/VX74/uekr1HOvOajYCAQBqhDdYCJR4dGg
ajuuDdaK/2zmLVL+O8pmXNs2OsA0WqGS34X+esSazHvWUlPrhV/Q6d/Fz6fMl1CBgcGUpSUt7q2c
zUCO9Qe27iK2ZG3gQ6/JrZcSFMWMJySODVflGE0FGXYDD8Oo1/O/dMWQX9whpIvWr0/jJcBBufIr
vle0bX0wiIkDcXOox4KxXFPxSP4ENv7cKRSh8AyCTneldhCCgq1HEPt2kMmEFCQvM3qr5JW8WQ6M
1cJ2cB7y/okFR/SBsNZRSkha0mLqM37Nbu0+Y8A/dsQpnxXl+1VOKdjxdiUJthtcGdV9uacoaYqJ
lRgx3S7tHxPqxxJFaJ7U6LurYCpbCGgVEB0hOJUEHYn7nHGsvf1UbaypUW0WioJs66fKeTyw6VI4
sm7TQPKPzEB2kD4LviFDcIL9fzJ0xNez81mQKbNifisuv072Nriq44xCMR0BWuioGd8ecgtwc0jo
uwQEdF04PJImMKRt5QlVTBf0RG59DKb8+cSCECm7UspSOMvTmokaeVoetlX6m1BPIIXjezdTBha7
41Ar/U8p3nW6dEofZDznyF1s7WVzKLvOonZilmgAeHNc2JEePV2cWcx70xfz/2lyH0eU9kBg8npC
389BjrIvNsL0+4gol6FA8MK7SlffPvUxjC5E9t6bKXrYBZjtn0qS9cidU6MpDaUPxKtKqndCzxi9
EErcj2+vdoXznMeODX6tBDN6Mne9dicYuiZ3lV0chXH4fr5XXvZppDWNsV445P150/YKYCFR1U5u
toexXyaMdxKMClXNYcXyCdbavj0QYq23b7BYdz5NE7ZKetUUP9HqSpcWCpXPf202OaoDIgOTu9Kw
wAXU5tyrphHi5NfMheaOrEK/C0HSp42YLZogwjKeOk6mjcuJ737gPRGzgUIwdBgR3cVSbEwh0Ri7
E48RVoxTYkXwKfUPagdCem1hvuttC+8uccu9UWSQpdJ4Qob1CE8pXDJUsPghGyNWOomdymViuRg4
WP54NDUHsb74eIiFvaK7eQOPEUlWzZcPoO1mrDIws4DOUm5LXjBNFExQwCkY+o8yt3i6dfm4jiAZ
pD/8vXuQG040hNLtD9Lj8UekdghOyyuqQHi81fT0BmHMqUxGJ27FZntYKJzJlVVrnyGdGrSBWfNk
+0hZnFRpglGkVrS1oMT2Ec3zlsea5i0Z2utyANoqaJnfAMBHnu5fa4x3LvT6CXpLH8zEfMB5qyYu
TVUVrt2leoJSbAsnhlXRb8qwgY8poMuFVFQoiSrF+s3E79+Gkf0XWJacV3/RobMPJqVVCCkR11+S
71Fmka/TTFUSx2q3X9uE0uEs98R/ZD7KCVWaybtXIxk2YxEV++ag8jNfse0ekGLfEIxeyVmesYZ7
PeAxSIswQAg+MwYZBtLLQ0cYXJUEAEDGmSFQ725mzuXcUsdE9HqpBNNJeSaF1TZQ+99XMAzRfCbg
HeD9DlDwCCTauKfIaC3sXgGObo5zwB1qApFnKCqhh0tptO19bhJbDdU0Xv7OBupZPkDUDj9dKPxT
SeSnApwY8N1HybUTZA68VOwx9lhjXX2/n5ae/pUlsLd5P1EOn2a62R0rprUG1Y/e3Ngv0pP1r24u
3iWvXaBoA3XKML9Bd+wFurI9YJJfoku50CTq26DEJluZjpECv4DKuuvupc0Cz42aXq2rFOfJMbz1
Y9vHI74UdRTuyBoCE6d6qGtlBJlYLd6YKqmkqfHjSlBBAAfU2bH9sI871rSn0px+KSSD1/HShStq
JgZiaw4JtiFbxJ3E3v0yoT3yIXngkHfLyHVEHhC8kDdl1Kn9YsIG1P6iUWbr631AWibValqKejmS
184uWU8GOQMu7h7dUN2yTWlFdzMi5UTAmdZEjXgFk2IftPAU+esfkiP6JaqsdyT3xHtKAPQSnR6h
HzDw8+UmOB+UxB+pVINHXOtiuRSSWBLNVSZpZDaeWDs2pSdBL/RSmqCOCS6SpQYgoldF0OjyIxRH
N0GPUyjyMyOcNKluBWvirioATejrigDa6PYB7e8IzLxGERQOqOgBPwtLngEzkI2zpQsOm4xeeKcC
wHD/sL2y/XVkLSbaVrgsTQxgEgzT2kycAeZDbf5+XapaMClIaDeXq9Z6mlakoSgSoRppSSYGt4F4
yRd0xRKBcO8WP0W0fQRPcVW77m9n01x6VRWU/IA2Pd1FiH0QCP30NgcewEYyyULPOa101gFJNelX
k2cOl5jaXB/EyF4Gl1fjhaAQBxe7mz70F76Vx5Ke2DcnDSrBL8xSwQkOtGj+KhwU/N+FcsfgV5/h
RHvRGiZe/SArN7H68eQsohocx91dnsjEL3SRm/+BWOqo4G34kNbBuiI5hZxZ7xNClRp3S340cqjo
s8+g+Shb+xNqPQm/XQKEBPQ46eli1gjt6cKhn8otSIyAbLwgj7kOcYWBfl8vZT+IDnzfUAuHauRY
qBthFU9fue72OEBESWgMupDXNKdUb9eSFkvmNRHHRFc+l+sK6HAqNREcyt18yqVPestFCLXL+37g
0PIAswijZ0de01nZHDoNtv1/lu8/bdZxhRWj89MPtWWiADcf6z+/uoZiXtBUTB8OkUcTP04FNx9s
IXYxwbBD3oyNIaszmTcn4zoa+EzaKGF4kZryKCurLbl5vJDPHOgsrd2uwXNkQmekPVbuBkx4DSmv
FvAb9cBHacw9zxgADPCrWlLg6nxaJNLUxCr3DnhQSybPFJuzrNpm+l+Gdy5SMsxWcFCA0cZOJgKE
ieObVTvhCQkZGAzU+KujUfWmhsm6oaKtAJBdRgIpoE/4lFgzA4FmrLYndkL+dmpYqj6uuGuzCbgd
JoTcUSV2oBc2lJASEXQcdQuCv7KrOfzwUuPowbujZpVlSUfzEEU7SwgdcjmZLhzqLSYHx2qCoS0F
JvjaqpCSqP1lq1OOJ+J4F3L9Ipmwvh5vmpkK15zEqtPV3yr9jByWwRoeiCKnBZPbw1rU82QliKjr
2oGJC0dtKfE57uO4a7IPPh/x7NDdbp8US4qLm+r+icYvZBLPEdQwGF9BpeOQ1n2R4ur+SWsOHCZc
SiDcXmI8pOEJ7yAnKGhsf+jmWLDoIT8w0S4X70nRtUZ6Zaz9fL8SHZpljLZ6yP0XbdMZxwru0Bdw
VvcA/IiWyq6psn4xFtycIlQGHO1BwKEguFEPKA3AkGVNG/Hei/k4P0f6Ghp86BKBgCkiMEzNE9w1
mFZv6l0XvqlUt0F6VsCgtJcDBewHCCL/wet5Z0iMThaT1FqNKjsYNhglwwUekSKGT0U9+Zaf2/BY
fGfkRU5jaDxNDmL9qUfFlQXhJSMFhqWTn+iU2F3EkDqmXz/qfw8UKB02AjHLAjAVaHufxeZ6zGNt
y40aNS+sLhDwltAC5amrjs5Eeu6dnbI8alO/JvafU6XnzwOj/OVLn6Qz1RGA0e45XtIGDhrcB+9N
+PbAKvEu976FZBJqkxpLiE/Bugwi9DI9MivTnMTqVR37EdDTdhFPWDdaReCYjiI/mnWlmtejH94e
vFones8EoEBRIY99zwZVrzcbrRa94lz/Y2wKvqu1QDOQqbEQYhWptyXccomZUXPGmowS4+aeauaT
IGHRQM/qEXmPMw5wVNq9Tgc2PX1yxKwFUQhRAk3Uq7LFtw2FE63gceZfdT18IIg8PoR1Ib1lR0RB
iFclbH2K758SG0CkPe+Xxxnr6jICr6lsGKHMpv2iwGgEAMha5MuWQqN1WQq7VQtQe4bfHhww6+7k
+gXDOhGjDchkTAoY+OJgcaJkip4tJHFsMoiA5rwuYhFZGptbz0MxSWhwpcl6m6WXZk5LVS6zDLUm
uJiUUU1EWTeCPMxAzojItNdZy2gaxnbfIaw98qhgGkByDQSXxhqoTnjk9IfAvhK2TWAMQlQZdCY9
nJxgldwC6YwBacEpa1J42If5hKg9hXarIowk3LEpQUiL9VKBo62pgXVfFnvfOrZ6SDA9zBWA4rkF
sxjTPP9zQrl1JF6zxi85I6OTMyztE2+MtLVPXTjMd+ykDT7BJQID8s2qUYFGY+TzQbD/nzW5D8PZ
TfRzJC9IM3szK1QIe6L3bJ56lhT+k2sgG2USiafBAE4cO0VPBaid8U9q8uOgf81VY85ebHSK951T
yAwg7q28CcqxfqDUKehw8zn11NLrIheqXa27PvcH4RadfBKOt7B2e1cbzKBr8rpu4MH1KE/vrCUu
U4De6rzbbBhTTEAaS4Bb1NSyy43KaOyjTPZqyVXRYt4eNaFkSdL313XTlbS9Pgtz+LX1JgTTqEs/
XUay5WBJReClHQpgBa+wgtw2CNYCzMQotiN35TtcwXz3wPuLj9FYGFchq/ESWw1Oj1KrIBEsJznf
yzbZQYdQfTy9QjFYpYjWpKqw2lYaM4vBjqdQLczGkzgEddq542GMVybvY7Zf60kSSishLncgAhYF
T3tq2TQwbzEnNJa+fu/jeT0sfNmw8dsv3/jupHMi1+OdTpNeDwyiwhZ7uLPROICsLP8+6x80KSvH
QmgA6X4kCD5FwRbCN5gfnsyxzX5mVLJM7eCrubOwflSar0X4gQHQdsSsRNOpJEn/3N7kp96ZJUTv
Ou819+sygQOO8XfLZX9Gb1+vycCECbHdLDTRf9Jov9dGWtpZE4AlOB+lJx93+XvKylXW7Ep2RkBd
4QZhZoSAGPv9kUASFciNGGVToMXQOLIE/3rFD4dDV2SJbJYEkxSpExssv52O4PvBLWcQSRahWdrd
o94EhtX+IDRl555ICdiR2saG/w+KbHzNmOabVT+QheJZg/zjEVFCJpG1s+JzXVDWrjs6Bk6XGEgL
uho6VFAbqUBQzJl/IQLTrQDe4Wg6a+a+jdv9WM93KSBxgHtKDdnGc6fO+62XSxPf5L5qBsHfvjs6
7BIydwZnoWAXABzCPfZvkN+Es4JSyF0nx6nJeGEcGg1ZQj2mJiDtGKtEV3mIK4TR+8wWOdB69rD0
688378yAyoGSqGA41KwXZNEi1TjAVxIZAD9sNXHZdOiSIwOGsqzSzOS4tuxSiu+BdzE4DEDqsd+k
WeZrS4Tn+T7tPn0MMJFAHCWBjQYqIkxN9sOexG0BjJX2b+xEcsfMsKgJozuBgGBX0b4TLXs9r1Fx
3ETrmZmAT2YLA9l9QZe0tuMOoUmuBiFdHqvah9+k7sHVixJzXxFMBB7jKnuFubzcpbsZJCbXi+gj
H5WnRKf1gfnowV4WzjksHFQLqj9qUuGwL04FqUbNKOw1usl1MD9+ID8ohAQy3JwUSK8PviWWDDyn
VaIpTsLJgRojfxQL7Xem+fX6F5qqCwtygASbq320pumbR0OsiAr5yGNJXwyArZCefoExBF77cejc
vpDUvLDkijlqIriAEAN0JLGalq+yu+R8NVwJ4+uKNgDtlOoq78Bg/UXfPZlMAQGMCRqFqr1QCZgD
d+OGKs2a1rTESk1S8BBrtUdzT2OwFXUX+rjuTaULTnU9nCS4xRGsQ7+u/PxRl60Fk637sE+cbzVc
BL//89nYenWUajF60fmarXirjuFGQ2tT2zMTPBvftx6Gysd5GedvsqiAAIajpNMnJD3jzgSUgRrb
7pVWF7chKQB9BM8JOane2Dt6QJTcnUVrAyQOBWkvDzu23qloPL7LQXz6vbxtB5jxWoj4QzTolwXB
3/PbxT4rkUHVhAiwQEVojg1wJBVZXMH+iE27t6P8n6yEJfiXK/qVvRQ4mZbSoXXlG2QQM2hbGSDh
58uWimzy/njl3CGnX4oZvcXfthJksBdlbj43tKuEcZG16WwrbDvLbMoOnBm5vg/UPU0eCVqygG9A
1tlnpmL2oTGYD/ti7yKZkRGDODDAtwv0tg23F/T39dyW7djXV9QETd1y1kd1wJWjiPhoG1XrKGP3
EspbBCwZjWxNavGzpaE4ECNZSpUPx7jbxS9Umaqsa1UyYSrqWb503ba2bEe987vRU6kYWdCupSKe
rgzxLOAIQI2KyKM18Fpaaa2bM8TKC5tRyC8VLikVa5KwXz+QdlaC7Y6h86zTKPxqFlb69C/aQMS0
vn4/niXEhBtKhBP10KJGv21GcFNJeU5TtZDG6Dh3EQwAJC3vdytqLfPh3KCuhR23RiIxC8iC0x/5
KMODKjmAlhRCGh6NzIADB483c7Ab7xlcftWemXqHxZywmw3hJ/FhK3VZNNLyw9rgN8wxLLIXYkkK
UvcyXUgKtMk1xz9HdMM7kB9H+0IoXfijWKezT81cqotMYHEZ1ThFGJXaKX1tRVhNuboHZcd8BZCy
DU1Dg7YVZAf4NPv9E2Qc8BAPOuA7XT83RjyM8EIo6TrKv/StVJFkrFcSl2Gjv1VoLQtRunU++ezw
r8/IWhkYvS/17FW9f8HKB0LxUSh4EQb2XJut4nehpuSo7zlASyk/xjNbLqjFooOhTmY2LDwlyibo
794lESD6qieKv3t/fxEmXVBuE1EwWLFwK22ZpYGpgaAlL7kWOn4QyA9sKK/sLbKm1SPav1fFQXSe
zaDugJoQZNSqbmspXEGqb9S0oDvCixMv/F8L6wiYr4tMMrAusiZ+HRMYxOKGjTjnAmPDjKZ6ALNL
SInbTwJmiMijLMNwwz+H2mMOqA3e3H6dLnrDWcy/cbIvhKgCR5byVTZUTdjjaf8s7DI79hV6BFoG
hCu/19+8fFDLV6vVWSVRjH+7ArLlCdgsPa9JmOsK7871GLloafCJilZGSs34LAWJR7JOAgFlR/mw
e5AFFpeHlqT3KQYfBlf2V80yS4YrZQnEZtoCAw4eUhhbUSc2T0vrztGBB3dIg7PhHRb091M8W8rG
ZrPOmTPJSFLUFh9BoND49UfBvK0AeAnp0lXpRec6ZtC9jMlweBqZG9f+aH4eN+RGocyXLT2GMTdo
2ZTAiwzToVMRDtgTQuv9nfu5U6n2ZL0rRVVWJzYTFx1K60mRT3czQntfMCo7pFkFiXc67m4ME1zN
isR2xGMVAyaPlPXg31BnC9Tailz1IHJw/TvbaUM7KeCsXCkC5VwTfkiBkekjzE1ZFKoS9aU2fby/
69IB6YKvIF8aAbjQszqz7hd/eGW7Pz9RpOWwct7xQ/5fYbQUO4DqlQ0rjAvWwUPEkl34xguTltRm
1UEA5K/QtHdPTKJfaN5NgqQXeFU5L9F/mV+bUX/jojyooTWHThSA0OLVbnLMkjBRnYaAYy92zGxb
MsvQkvc0z48w8TsdIVjju5qWaWL4T6LnsooCCJWvv+i8EbL+LXTNOXAF5qF+X4DhDJ74awpFEt95
oFWJ+Z5ylDJypTLDLW1QXV4CHmYR54Os7vwTg/L9jaj2ylwqDlf/IXLTFlVRtTNzVJyUsaR7IDOO
KRWcWDp7OEPRJbyrJRkpuI++Oh7+qrXOZdysx95sZGrMHAQo5GJ+u0mABl5u4O/sV8Juv+cI07Jv
KEDyqf46TCXxIBBEEjqpNTNezgCXP8Bnsqv9scdKKFp4mXGV6UYmRwE0ZUTeo7djzhhjnY7EK7RW
zM03jcw4wO8j7e8qgq1K06XFhU+AS0yMdOtxBUkHmhRcuHNb6F8JC5/sHebK6Ar1SHMBwW2q4XDC
vR6Ss8Qf6RoyegLS2eRWTM7u9H1ToU4go0P+RCZ0y6RZAT8VclJ5P16xpxwH7fDef24Vp6rQ5mUq
tlp1fMbmlrNDrhRlBjIjFYFNH69mrJIUtIGCoy7Wb3e94V2aF07WSwzj7MNq0ZbXPQQ71YKBk5TJ
Cy9smGhUl4GCDElkk1E0HY8CTEVDq4y2WvvkHMqjfmPE41o4smltQ6omE8L7HvTMOZ+5tTeKeX0X
r7niBIKdg0f/C0WHEEULVGsVWMQl/dHNTu/TUylXuigc+Zd4kcMEuUiKSBd/hLzfwFBdmyERpD9f
+UJc89j2lXglQJ52qUEHH/THb4tFVMFQjUXLYu8OfqEZl6XBoGnujI7XMH9To/hXwkdTwtAjz38s
fFG/XuhJ9HRUNYKyrhVFLKc4TkunXJ7qhLsYe18LwDwSg4W6OyGcn5kn0AxVcAYUtBXwLfMC8QfD
5NuWdlOg3bSFPTM3NoDg9KNPQk/Ov5a2khM/1xyLojeuRbRH9vUK54dYx0eAaijXKSrz2Hd1Gbpb
Sh0fQnIVeUBAR42i7sft2gkhZd1baE4CwZD7TdUJQVEY5MqzjXgD+gEYN7hBZUP2TI4peg4zvaMk
WwXtY3sOF7XDze0nyrqnOFzeKXpGKG58K9Lx2jlGIkN6tEjWOYz6NzoxUljZcdthV3RHDu6P7sSN
BpckJ1JUsE/nrMy2H3W3j7JNSPeqFScizJ8Dzh1VGcbDM3gSbkNIUy9//eisTsxWKbliHlxXyQjx
lpIoYLYQV0/AB8nnq6R52qyWpU62hn7Ikk33eNExPlfCNB3co2cpxdfkffYaS4x6q0PF0CtFg8dZ
KIWb5yBMnDaLYnR8O024zLiSSJWwsoamKK7blYiGMbuR6RYWksLLNmzVhEtw1925spIjydCE6mOo
V6I2x2FvWbxyCl/pzG1zDZ/F3XsB1keMqzHDeIygG2VL9XF72f3o0xltLY0uLFdkxJ7JQMxXVcvT
YljCrrrvLptb8+fyFnW4PfLlRKQbX0rt5ORFVay7RytqfPhr3GDJFNGmk//c8yIojBS31jkcyzlr
dhSZMCPF7UHg2v5ZiV0EX+G+vhgvJF5itDNhhMYo9TnoAuiUMUFDrKhxa7imkL3yiEUt3pIdiMUD
lb+3j9Tp9FQ8flW+DV7tmx6AIqv7KCyI4f8pVedT2XU78Nc8gEzX08Bau1yvwt4c6UHaHVDjUdAC
buS2bgicRaRv3hV13gaVsVZQkhnXSQcWR20qKMKg4EnfO0z0tzpbbSV/i5trSZkO7bejqtR0OTSz
heXZm5ltYeGWl0nmyDsi7wfVy55pMfg0Ep4mqmAzcyjF8yDRN7leSizrMsKbV6y9l5Yaxb0e1bc0
/cE/Ktsx/KHiE9vafr7VeKK7OsGenkmgqDMFrm9JZDmK5ksI6hhOCwMKJ9QZAPP6Ch6oFGcnYpPt
JaZGITvxftVgqQvm0Wpkly1OdhTsQTfnzDflCEYtWl+Y+caM//k3xLUPkvhrrERADrJ/CkLNExLe
FVgjbNl3lnbH3qRCFwQjztd8PW7Rn6pWp/iaBS3Ovru0c5Tfv0Li8Y/QDsaIRd2jR7pad1PHBByd
Is/GUKuFBkbhOgqZKURA9WLn00JGgto1XNQ3OHBQLfW3nGjJFgia36OBL9DxCqyWx1wBj28dsIZS
oTnlNrJHW0+GMEuAXrXSnrqPZuFI80636HZnYSC5X6TInCM5ZZs4j505ZnNLt5NEnjNznidBvkgV
0oRLpJJi7K8I2DniD5RdhJoRE7u1tR+xIqLvRthfazgoKVHyq90IkxXq+cMabSXXeiwDE7tuW2Yj
hYR34j6uxGIX71Gh1bT10MCvTImjUPPO9fgfpcTx53Ln9BCTDLSGPkghXJgeBN3qog26AO513xp+
GHn+a52f6AQMbZdcLyXfigW+6YTo+SvB53hdv1WCXBQFAlHewYwJ2zzy2Gg8CRzjzIQJg2Q/rvG9
C4GNLAGLpKPwKOCEusnXsbZl7R0V6zop9VfpvON3DNMObmPv4DBf8J+Rca97Bj8gOcGkcDmsCK2w
bP1B8ZMR+NII8OiqOcXDIiiew0w92RaR2CIu0rM2+tQQESc6D//uwNEKPOB+9VgQ/9R8WL8gcNK1
PJLvGVb5tVKgIRVN+N72vbneGWwzFeuU56t1cSN6wWlui0mKA83D3QAOOBhQYVJlapRHkZ36ixei
ZApCpXVOew7X1crS/GxVMPtlJzlhjImGYQZnokj3LefoLia4YN84lT1tSP2uifIH90qONj+XC9Yj
euh4A+2IpPqGIzNtYuhtivAdjVxCEP9lOavIVwDrKZwIvtUbkWje4qhgQCOK1eg+4LMzQh1DPrJk
S1I3eJRoMCIj6EJVxMYyHcZuAg6dUf1h268jNlNe6m9PeEdtGbOWPEBeOHGXZ1N1B8elXteuRLhF
yv88VHxB11TXV4HJN9RVxg0QRBIfXOdeJL7j/TkCHJMq3ZYKDJTLGLr7QE6S8cV+ImEa7D4IFN99
sQreWTGdKxaZ/6groKmBTa/I5cP1sbEwoRJc9KBIY1X1pQYsM786eJYZcQcLjC4y9S6FysSBVZmH
CAg+SjqPRvtpX+BBKeh7bKYc58yKXjN8U69KZYGJMY79ENLcIVyDrpKnnFsZh9jUZ2P6Z20Z04W0
MlkE7u1oTw02kUHWlmqq42rTMWlZV8Ll3Y+kJI7vAb56Ejdqgg/3/2fg4xH+tz27QIchbRpF1srO
UtmsXRyHtLtQ37UjKcNenph0KGiacjrczw0JlJR5QAPR2VAg97qfsvGF9Ve0AhcjNzjltJwYR4f4
d7HTOtYG/mH2VP6bc5bUn70Oufov/+0fxuk5FFeF4LUElyBKRvuYYr4Pk8oMtSikbiw7ELNNGrlA
E6G5WKV12Moj5QtkRaurOFaLy6j0eJHtEfs8g0ULpNz0JaUjAApxrzgoIwBVAcdZQGQ6y9VtiCze
fQiPKzB+gczaPWOu49VP3n15KTgjJwVIOXKr1mvSMdQkgGUXbma2VrMcmAo5wFhRq8WFR0Dsi/Wg
FAnlvQlXbQ23qAwF2vEq5vLhBVtScpS/UNIZVWXfLLX8nIEXZYcSyLndx8WVv0crWaFAW9hoUbsN
T1BpSMJQmvSd3ycASgTW2u0mEk5HZJb1VRAGMtlPxq3LP54N1QkzzlJHTOchJHZUKKX2uk/nHlMD
N7rtAWOQJCF/U4AJHLe06WZ4iTZYpWfRtsP3Yo5479gqToGPXECUfVTxCPIQgKPyTrYKmhhzreLu
87nfbC4Cn3LROKAw555YuSLdyouPUl1uXlcfv1NPh/O2dPPTFmwLP8sKOhFjdDNv3u/wwhjodNCw
58xR5whjI+3X5/76cyYbQ5pL36fkmhNgE2vho3u/+C3K8sCjnDnR+9ajI0zqHQpfneR4cTemwOPn
KT+oA4whOigl10OvUfo56arakzf6WqQbZUBeHbhsuZO8RnhMwb7Irb7HCfh8FVJOqhBwSLPpgF+C
5bKVaQ0goat/TSIegpI2wVyG60maRWzOkpHun8nvSM97+PFzzBelzFP3Rk0m3F8H+nfWHWAvApdO
03KCwQRP9zNK+nnu4aJ+O6z0r//wvrciYZeEou2j8O39YY4PQ8r5eQnM+DUVk8Sd+Gtnv9V027Qw
GAK7UviE9u1XS6id6ilLETikMUf6vSONM0SaXiEXYVXG5yHVZ4Dl0/4WXrrS6X6K9tny+Y0rcyWj
krcpyD8FGrWpJA0X5yMp6zSLB7MKD4uhx3WZjQLLfkYxTXh8zt1GONO724N8i9H/Ss1Ygj4g7Cg0
XtsbU+dVgk04eTcQ5HOKIuhq+Hv+9plheGtapWGErctPLrT7KzWPOU6DX5ggCV7uk034L1IlkbK8
vhGsD2a/6Ch5XBP3+TkCz5eBHAU0RDjYkLn1Ba45cG5I2mKMJzTm+kpioLIprLqk4jLgicn4WfF/
cYTxfIdutKhybyjY0obuISsCCxG5VXdBUrVOAFIdGuAJLrIRouFl6wbwEkJhgFsTsyaixslDA/O1
DZea9NWXwrFHBKdRqmFL23/pB0cUmcSpTZnXJWZm1kDlYiZcRbhPi9FWcdLzfwMoE1AmBIsxlh0f
xjTwRRAdb5RMDs20u/4LvrquylWTeKTR4vmPqA1R/VTi5cOtCTpZ6e+u5KvrdCGkIzAh5kHi6uk9
8zknt1xA3d85E4xQoAsJPJKA0q21R7S88PD9FsQFKucM+reFy71KTyzE5Hthjx807dcGe/KJYHF3
g87mS2OJ6GBezxmbIzhRuFjfuafenaIDS5yDLpoy3NjVUc70wIlAKAol1djpvAFJu3M/S3/6pcpx
7nOXql+wR6AuF+Cj1spO6JxNTN/gBkcaiFqUZHtLCzog1NHnYKpKrqRT6w8X36GbUE+9Likh3CGJ
LB5GNppoEZInk32CDzGR6/xsrXAVIbJiRWwHz9jCeNku5oscYaPWefO0UBkGO7QsU9ujUnSBicKp
LfFU9sdVoNbqe6az+V7vW8cHim6fLnXLoZWyiETaDO3znaRtb9m+n8I0/N+ey701gAmwQpW3yhvl
LUq3EtdwPlW3cOlhkt/CgfHICGG2i+J5QWh1ruPg15uwQ7Eh1hSm76714tF+aBLw+LoyK05JflL8
1cmBDJWAQr7qi+5EfN9a9rSlFvis+LTIa85Ia3dtBWQgpZAfndCOZy+m0nNcl6jpv9lYDEQXCa/C
iv7rYMvv7xL7YI0F75vZ986vdSvTTTGW2aaPYuM/Xp2bLMgJjiNedjPX8L6xxB+thQFHnSgOdIxi
kvK3bXzJaJqR4UQiqNSlI0B2FcCMpwVHuUpjldKWZO8CwtNJVAFss9spqs3BPxKvTVHDnGDrLilc
b/ZYQqdrOTHaCUyvH9DViBrGUsMh3pG8LV79CCwdEW5gKFeIn3OxtMBmZZtRtHCzcvygEBRHwZqX
4zQSnGeUwtHXsehwB4gMFl0ivwtIh/JU31UULzO8C6adU03N4ldtfQlo0rbJXZurKECrxszNkoIf
kXNUPuQRBmU6Nw/tHfwFfWviDgCg1bL6Jg7pzopYCuFi1ljlEmm59dcY7ZTZKhRcTQeQTKxVVg+X
IX7gymrJEvqZ4MZ/tLTEMAZWLU7pO4yMcDVtxLn7AEIHUSOkJQmrNwmNTC4VXllFpAiOCQpQY2Im
Pi4OvXsTi9LMngoJvPOkQQrMRSqqV5EaSiSNeTa/q7ZSD/gkerRNcDN4hMq5kUmCyD28X7acU127
O3ATNQ5/LB0NrCz1zJyEj/irr29QATaiStWUlZm8mu1NrIZjplE1+RRz3wE53qn2GhEm77BO7L5g
cKZjlTCoQW8Hhs0pHt8jwjlpONL5hMHxqb3v9cZA/WYHZxq0lP7iQ91kICi7UxyUyxXXDBOgRbo/
h1kWuslAU8i/2pZ+9RbeVsvrZGtvCdAGTiZU2omL4G2WPs++2rYEUsj/dNYrHx90VURfYgXE826N
mzzoDPYWBHSctaDbu4X3uJvtF3b20RavieOzErdqB9aDHzBN8N3OVjt1EzQO83WumtN9vYN75WGp
9UvARxdAUYIJuDhHEywUoALvsLdPa6v6grVOttT8Eqk/BWe4nOMIoFOUyRnyfH47Z/iCQJwxqxpJ
r2ICkIKz8TkwqfifSSjSRPBZLsAjAc8egNrOxyOFEDOIJD+vNLjDXYxwrS42m040ZRuPgUtAqrGq
tUraeX7Slybpiy9PdLLf7CnE7Z46oZ0l0r3YO1Hg1eJCE1LkzZT4cKfIaxcQwQxvawgVndEoSriF
pUqLM/2PTripbea7Wkb9ULjnrac+eGQYPTcGwib9g/08xeZmiRVIqXkYdZ8Qpq8PLFo44x5zbv09
CRzbp7vQIZlS4T33TfKvzBXmEmeQ3lmLoNqeXx/xP0p482Lb4UpYh8E+3BMSaFUf9/uenzR8sp8N
aLhJ+FsyNa7kplD7Yw9DyTMaUW/784RYCrdb5EhaRvUTFwKADwBAF9GQimpoBtstLI0UK0Bj/rL+
sai1IAYGKudNBhI5k95cAJGkBw1PDG6R/IK5oE1Anj3JXswum7kxTuTn6/uP+WYW0nTWwQ9SXFAY
oCbX1GuFf2ByZxBsnFGlTrN/5EdMN8MnFVeMQ86BGlN6fqOKLV0h1zTpJq9HOGxYNp8UucAzLxrs
Wcfjo/IIEri1rRsehpqSjnVMVNSnp9toxKI5BHPs6xj3afCxob6xgioDKiQaEAMjjJ7gTWGZH/8Y
dWJGgD4uMGa1wO0Is0P396x2xbod7dqom1TPxMvjBDa31h0/k4EKi1aPtPCjo3D0sAxLcFJyAtG3
vTC3Ln+d/Som7ldWuzU/abcujU+safJI6pnewGS/Jv3QJab6ebLQsN9BcE/H/DP+B4wECk6LO1Qm
0sjlhNGRy5WDKAnqwZgWm+ZRtmRP3aTvw1HqFdX/3biqmAzqVlDI3An0ex4QU2icd4QaD5Yq/quW
382Oi7zeEU2I6PMiBXBrJDEvg4JzZ8M6srtj3jneO7Yt3hXH/7njtykAeWe4kcjRqO5rOM2k45Rs
E/lirti5vE4ow9PUkMICiNHBNF/N4T78Uw2uMIGlM5FMcC3g5e8YfwwfXqQJk5ayylkVtY0TXYmp
hhn0WITlhfatZgGJH75aqtRkjc0JLa0bya8LvseGf5ApNzBTqW47RhJkfPbdeM3U2/TpR3TF/ZXp
tvIOVRGCWxhGcRR07b3FvliJTOKO9/wjYrJ6K8NE4MaFeH7b4PbcPvSeTW5BAiAdBkz4+JkawWe5
7YSqO5Lgtkyurm2zBmz02zf+5OjbIEf6WnX7B/cbzJRwLSe01zwqWFh/o6+cHFLbeV8TMg04LfUb
Ar2a1w6DnLYVzrBuvVVHr0/GIVMChaCjPH8HBQnPrKarpZ/ssC0JPARRtGfUN5Jh83z/1l3d/6uj
BN3Q60vZjMhqP8BFRJBFr7qsep/+9EkLuqD2KpYOpxlxqPE/0d/HdRACg9l9VFsI+NOOVNTGjTEy
Yzyoy7hegU2keOogmVvAL1X5HMOf2OC6d7bR8lEtSggm4zBJ9od0NdJgtvlKFlcnr4ZyaEoRx0Xg
HrgPAmgyivd8D6CjrRlPAIL9oY5BWDxH0UO3c97ePPbAPaljCHDYhaALkqOUG4jTqa7yGrtYrTE4
Fv323SI/b0x7XPPD3wu6qSsHQsO1sTVr2VfhiZoHTPD9aOaphq1VL0dWknclYwvpdq2DginXmKqg
qhdInDysyiOrVEDy+BmyDjgD6q03+ZgGhu7R31/G07EhEpNZIVuXBpnLYROx4u7GvPZnbf9h70ZD
AAFmnyK+z9Ks+XnZHZlA3KXTOHe/Kvdw62CT2J6Y6eRP9KdltXbmV6HXTUXkjUPPrlek42xbQPrd
JoLLR1VGTdjaVuYr/9CPrq57Tasac7yQiNp0kS0c/AcTrGMZroHo7e7Cvvv7gxFLGrFE/B66Kzu+
liozQez9l6oN83r6hWILPgt3PPymOSkWRUQ5Ldb9HadEPaC0YmafQkLCs+p4k1uU3l3ORFm5cJKE
s4SHKWIG4gQDRBsydMlVbR5Tjk+/dfnJnFSOzLkLPYU1NDwXxanrmOFdr+1qkhG+1FUkhaG4icjA
Hk75isL6ragGnig+E8hixOi742Q+9Y2OyazhX5/6quWDd8VOiCsfE0IlEyQo9XJsArft4HaTOika
DcCikXLFm/t2h9d2k4axZpQglsO2l0EF5P0/IP1vlSIR3LkVQdzImbanCRCa2Thu88NVPNLQc9Ld
jPOjiGhMZiLK8AQvQA1EgVtnttc1jQNuqGNUsP775pOcPR1S85LkxM2T+rsvo3iu6vAW96yGHX1H
raKPKb11RMElL+8InbYw3GsnxK63Dbdmetm4oTtYyj0prIiquK822rwF0sYgF0yBmYuewIVFnLrC
HeDjsrnw52da2jjLg6OlavOY5CfLYtl5ZHrYOqL0FnY98UGA91snpvvbPF8XfuYKJpfvBU7u3yxX
Xt/W7ixxs8tafv6KL3pts+0lqHReefGcKi8q41lGdbPsbfQZwJdF2z3QQDVi6JdrblD0Q/dT+g9L
FSgiDiokYHmy92jn40ZKQSpK52PmeJ6eEy61IV/f1DWV0efKXw9FEM7jMkpamz49Pq3NxoHzlwtn
1YMw5hVZx/onI159SrVnto784FzNGL23phMu0rgvgFyIh3RfDhji6bkdp+3A9XTCbIHGAbsezokd
RaIRHqrhIooOSS3v1N0Y3c4tTspMY++Btz6F6LWWi/D/Sc8s8JWBlIe1vOGPL+xw8fN52fXJI82t
tys+lDg0fq5GOCbf5NCOnVt9ODjVd3zb7myQcgjn455UACD54C+UOhEWMmiQWxNII2l9tyl1QP0T
tHsokwCFgF3hFg4KEFmkQC2bChascEfkJzYZ/I7rn9XvjdUH3GvOa8vq6ijb01vPpgYmFaPEZ/hD
mMQPO88qHIA4fcArICio/VAjO8NGDKJz6znsgKAEM2/as+2c4KuC9aFPjBG2Ul+Ur+v+ltM4qfKN
uIwgsF7H96lnuemaaSaEpVUBWyf8tx9JAkBnus1Qs85Iq5w4AK86hvQej1wU4a0ex6uFFi3lJkGj
ZnSqbZ95z9g1nd2ns4wHB1cTKL8PX73p1uiKN60fyUHnaRDtt7SoEIm3KKktN6jYSJa9q9+/itgJ
W/acwGlDX4/mPKOJNWR84qeKM6wuoGqF4hhBHzbE5rxqtIJI/2KSgYhuYYyfTRcYKAUnN1Rds3Vj
uvfeznSVo2fUO6pWIKdF6zRL0Kmz0CtDF169/kgWJNHDHwvhRUVuYXqjZPCrZ29BQ2Rd66aZGhag
fOzvPhrfESGcWd1gYn5078Bi34N9FTuZbbaVNgPCyQB8MAJH0yqfjeEgWD/wMC1UQY5pmDefjEai
GfTjeliRi+6l+mbr+oAmDuIUo7QD8J7vaCMo4CtSSKLLHpiGrDW9QTGHhVbxjIE7HMVwrXFkzMwX
ONvZ/TsV6azrIf6+9D+ZOcVrFGKL8gyz4IcOrW3cvYOXtQ6grK3oSprblkchvK12HH7Qkh1qG/1Y
YkE8bjCoMtTvfR61L/OgOhOBjFIy7jAvKqpQJJ5fJU0mnb4dW32e1vDrkz+2ag59pZYYrOK4S2k6
zh/x/7eBv9keb5RuH0HmQVY7NChCmxeIa9pZZGAkBvGGo2mw/bCP5T2kk/AMJ2+ZFKJx5VnZP7d0
TNJItMeTUp8n9/kV9GJCu9/npYekgtlsBtL2gCu68L4EulrZaWLNHB6YhI3BdJeKu8Lw6TFKkXoe
eLFLG2Wf2ypb6A24g7euL6zrCTMxpo1t54uXL+AJOEKMVnVYCC2yax08rsalpvtn785/6hSy4ssj
bs0oy7Bjx5PEf7bZa090iriRG7VT+5vrZUyeWnLwAYlnmoVPhIRExB9pAuBB8gQor8mZX9hfgLoj
j+4Fiwsx46FmaaEQ5DP+E4EF37y5x6sZNKV2WlW7w6d+LD5q7AJkVppX9d89VTG7mH/3Y8IWo+0S
SvctFNaLcDwBVVZQ6IZa4iSI+xKkFb6xWM7BimDMXMzR35+4d4l4CZ3kmzAm+YfxbSlE/VHktZPg
QQuDdU0Q+5X3rofvkJaN1eNFIFsUg2hk/t9cLKp62dYGc7fqpeFYKX2YOEm1HQJntmfrMwsQtTq+
7vdTE3j3b4nqD4dNpes68igiTMpAs+yGn3u/bEkjdQgivL0WkkWRCjgtpd2H/vSqC44FH+RGhRst
6ppq8V4JMVejjRUvt6NV5Kh4HGgW1yaY9zJ7ZxXLSuovPC75sNrbs+0sMkt6+Z3YDJwfEFXq43Rq
7QNyoJH9GY2DKJq1dlFtOqM5OdYqZzROaVPmuzHSXIs284AgbH3a7T7XgfAf/6bUnFnh5WBS51lY
C+dQ7V3JJKnjRZQ3HtRi//ep8mdEAlT82F5+d27R4iSB4dIkoePpDLLBi73azhZ8BAppXfn4P9JH
Zl5t3LFYlt3LtBJ7HMNjTSln5grzmtcIHaCIokXRMLY6FXVz7ejRYlFtR9J4FHCneQ78h++OXO4f
9Ejh67eir5ciXEdi6/A2VHakIMDkRKKK4hSehWnfkQN5upgpSyeeC3UUvjMGoxWxFH3RMq1hToiW
qnFlI1L9jhOEx9g2LI0QvkfT6fL50P6p5xHlcaRTPBzi2UbyS43eylGc/L8zFw5527zTQDtjKJOc
UmaQV9bvCMU7RsHm/CeyuP496YE9gZ1xXAa+p88A0Fwh3qHJ88O5a8R+Ft9q0V5mUfoc3OpDVciS
O+sin2WQZtURjcqINJfWHCf868cs9n6rnY/bI9VcIEkDnmp8UCJ5zE5UR6PBV3D/Fvr2IZfoYkVQ
ad9oaBiMrHbtmoiP9dzPtiqrGbnpDpBxE+OFXRw0VfhiuM7Od5rh+9QAXfqrkAYc51GaDpNSn8Ub
uFGlRGbTBNhTnBa1GdJqMtOvcwwQvwRzuids7tk0IyLmZgySVSfaCo3+utXVWsLx1xta2j7Z8Pma
RtKF5iusdvEVBzk1uvLRwJrO6+ISVItRcCxYKi9SltphwT+6jH6vvLt9xuMnzAvD2UpRm3fHbElM
2f4+9ppmLGzCZ6XkXf9h63u+LHxL15M3aOAnpmdV8Ngj9z5LnRJKlJbeHiJ6XV4cTfAvh79vAJWo
mFZUDWBIeUhWpSmD4mBUspUgP+6RBwh2WQENHuxb6W6yBAOxVdNvzjXMzZS9Z4cuRyjfSF7+CfPc
gbOGVIPXm4ZvrrU8e/ElY6Fjyb3hOgqd9Y2P33WszEvnhcGQB6m8x9LmPVfXXfBM5PIJPUMq0gFQ
iT8nUMfiDELBkrIjHd8K+XCWFx5PCPFltdCs+sH+xGFKjIYEcjH9g41BT6+98w0hEGnQm8sKwm9S
EPyUfvxLWppBIoPrm/eWAkcAVpGzTju3bAaJwBLBMQhYnuJGmHwAXDFsMmc4xGjBBEXUs92RMx3p
CSNHgfzNSLW6INSKFm4cOcuQOBnOrzjLRm3IWZ4VOLB/HigM9yakApn76k1uvVH73QRwhRR38rSx
pMP60zr9UgH4UhTO//4ZjdlFmRTorgKCJ2g7mDpYWX05bsHT4hrwXI4KhoE+cuRviwQYexx0jReH
w5vDv3aOmPUgsTjX7XSDMUzlsXZZv6IF0Rq20fLqcxP3OftKy8PfmMbPxZOI+Ee7xRMvvPOUNylO
LHhh7YTHkftXJNUY7KIdCQDzswXN/oaLOrSNetviiWYy3Prk3H/k7tGptRBeBzxdiLdzvjiBlWCo
evK5IN/0yISs5oMtDwapTJwkQLBnCKLE/itwB38LyhQ3mDycDEPx+bcQvB+5eYWkm2UiHMa4/M2M
Eg6fjax6PnoIY04We6L12+/BFiorDSlZkMg0MRqk+l7KCGeppfKR7vp79VFYaVEMNNW9MBU1r7g5
ImEwivkzkb6FPlKGlnPGOVD9mHp4bspL/a4B9nQkZ9rQyUmZVOte8srYV4ukquaSz0avkiYUThqa
RTJeNZhCPvYSQ3Bpo99OePWPSP6pBEUCInKUP3vsYjShVJ077ITCjRlPZojlWYEqZAz3aiPGJmaJ
YwkKTwl7SDXOzxBQKdYGI50F6tQO1JVIvrlFkJOcSd4qYs1FZppxqVufxhGxn6OwHiIgTT+Hn/6Y
V4uuySolYOpxLDRofM6Oqz5VDzWdZw1vPafKhLs6p7PGOP0VJfrkXG+10awSV/doW5aZ8qIcRlCw
UzYzxh0A8Bh8Oc9tMMbaBs86xSBMZzTuREmgQx/DURDpFCPShrH/kJkIc+Edst4vBlTzrlbf/CW0
oGT0V1YdtQT19ryAfoQtFRYV/om9WtoBBaMaoH390rXHfy+sm/t0G7UyxBBSvG34S7Bbmha3YuNA
rp5t81n2wrME//3H129P51Moq1im8saRwNz8BA7vNloBjkYG/QEWSEHGp+hnrwQxeQXYRv4f/Ful
Cwh4cin8smMGaE4PlK1x7mhDolg69D8HNxkOn7VPZMVUqS8vhUp1OmvWA+JtvpVUdg5pBLI4vFSl
kXhmwBgTvClZYIY18sBI1JoyLEqVS84uk1Hi5/+egiCueEkDYYrxNHtlSIOx3uGWdMaLdI5aEXa1
zr2hdXz3XbU83uwHI4zlVZF4Dt3ENjwLUt1w2JKthjoltYfFJUVy1/u4h+F5+8M047hrwRtsCLMo
KPn8WN+grAabBGJUWdUCwkfb0lwtvgSgZGu7u1YGYhkZ7MCAH3lWvWWaZD3ZvKb1sulkOHiYpys1
AxVHJqblMDspeebj/zTiOkcMcvKJx6P+lAOT3ngYSpL40OElHHCtwqI2wb2fvCMZTtzx42WFYTfa
6/6NW6IWacknsSqWCOGFZSviGGegcpuMIksrupi1UuVS548TygP3vZ59shE6x7GyZafHTMnFP1lB
EQbuVLFyJH3XwBIWbGsYIDkNvJUr5ugXPr9bFttSXTUXxmiNOYWDhJLe76EchgO/67zzJrmITJr/
45UOjeb7t8e8On6WnB97UjE+YNX2iGmHTuf7AMk1jxze4Nt5cUzRysZQ2LdnMe6iBmMl2U2YStnP
piUXZ5kVo5Vh1y3IOM1uGjVfpUaVy9QZXgsoZyU2JS/ubfFAhJ2fVdN+abH1tM6euVA5h5rZ2OWF
cQFImzvWiZXUc3AA7f2zv9fyCVhf/7byhMMjh63QNRjHXqM8D/zuWRXS0cKhedAovcHIWxDMwG7Z
0vim4wFvbumtpaFveq/VEIjqVqGkBYzAwSkp1GuxQvXPHVVMCn6sjNLKwukL4HW64JLA59nF5iWY
bAlL821bMJCqMjA6zDOtqmTgYso6OteJ5MzJVVI5etIy3D6pjQZw8tgqOzmaHT3D0XMH+C+IspwQ
rhGmEl5VmqHhjwUpva7gvPMyoR75B708rjf4juYSDuFKg0mCHPbsxrwrHcHySqqKuqMPfRSqh+Lv
aMMBS+jeavHCmS6p9au+hILkdygsuYkGSXbjvJ2LcIwuQmSksCkibIAY3rfcbYdxgqRDuLONdtpH
Falj9y8Hpa5vhypMx6HM3Wg5G6TnDYoeInqBh2UnyTPxxrWK7I/HE15YG8z2SnDZiYQRPcUcR0M4
Va0L/lv4kOQWLEjn4bRYmAhnIUISoJltmpX06ZhyOJrbrjkw6b8X7HqU1bJl9rQsauc+PlpJ+ieP
NLmehIa4snTl6oK+VQ/3ajlX5vPkvFUAncUdBxcXWneFyWDwtiOWQiWCsFM3mFi5lRZhBYB5dkH5
MJQLSJw1ZBe6INT3xDaK0i/7YViJw+rJpNxctNW17T8QCbj4BpCd1O5/ojYoJVmsbXJbyMPM9sbT
2RdpHixVQkQURS1wfn7mGmiONC+nH6tHnpyu/m2APIXmwrYFVscdtM+4V77EyTzq/aA6AyipH7T6
/RR+oIIf0WXDXt7fcFm2EDs9H8NSxW2XOTVe2ss1E7a08KLYYh9TeBlQN2pug7MRGTwcb4E8rD/K
U737sKtz7PoBuKzd/fezlR4yJuKZIiMk31diBbmw9d8vxCtbJClzPD8pm2s5JHHJ4mcn3DyxoTJ2
S1Ftpc2rVQtHEDMlxaIJIeaU3W8lRV1yyb30ZwlE+038aiwaLiUD+TPtgAvr3Fody5IPHRHTzWyq
UYlJ45cMhQwfDLk18bE2j8zevmVVArq/YSQd02M4Hv9PeHADShsmHFwFoXYqI72d8s/eikgqUeHi
wVWoB2JGaf7qWM9dqi4fvx734TZpOQzajc1On88u6mJrzFmf+mzMzGw8KSKg0QcKudJIjS7u7POG
nOeWuqBGgqcxK0AjEOLJEww+Lsh6vJt3Ou/kNWRIdCNfXyIvG7Zmm2p1oXXo/BIpkHYsXpL0ayPL
1BS8juGqfKLCWKSaCOm0E4Gu5k/uZoe6pQPmyNLMeVR6dCCR1pm/LdhvAaF33801pd0LfWpJ5395
/7TOKML/8D/M3oYIlJzwv4ZlWAD42SkZL7RE6FVzDk7RLVxQpcRh0zVW2t451bUdjAqy3lcV8etE
cpaV946nq5Twe23hAm1ZHl0V2CJ/UET3fBHgMqcaM8jX2prRLKWUtLbQpSJ3ZXrhchHfmSmSeWny
aATtpJdWlajqRM/BszL9kqe5cHJ7/dgPWsFLYr+fxm6UuQ8+GqU9qNXcyzbyYScLOaVdiHvUpMcU
qAuZHuhThQogtTMJb4yA3DNuumkH6tEzuhsmc67jvBRJOxBB3fWNmO3yPOuzH5Wdem5ONxjfUPHe
jiziZdmJ34HpgMTMrQh+SL0xCfEXqhOnCuQkpw5fxRntqbM+pGkJCMM88CkEgaVPhqHasZFAOxu5
HL87KTcp2IGjEEBZBRqwciIVHuKDcjxUr0lJB0UIMix88iWaVTcZZ0fYsSF9L8EyTKquBKL0ySWe
Lbpm6k4lfsPKx5lTlxTYQPlXxijN14IsFaJODzyfCBv5Dc56+pbFAR+JYHi+V+oCtBgfqk6a2HGG
6whhVy7gA1xERJgL/ulVVuDNUnoOrGdsLPJiTXwG/ODvhXmvN4PFhVigvFDX7CCim0ljAakb/F8d
Kp2On5m/aQqsS7jR371xqHbwty2WEkJraL+i3o1sZg1SGMOQO0O8aRQipUxriAebCyWiTpQGR6DX
AZHq66DVC73c0QMTc0w50gFMpbPEBVsNciTieri+QAZGsNwDxKDE3BD6EGTCe1kBO7H/4y6R+60z
GQxRKG9G4YWr+Zq7NZGiIWneb/hO8b+saLbjPjVQiKv2okThC1ecUydzyrcKpkQN1eOz93R5q1hL
p14Q4jtwbSTFF0UXpQE0qv+JrAnO7t7PT62Nf9gC0CPi7O5NK7pNV/g0Q8z6dTFsPbq2hBk00y0F
Augla+3IWIn4Sld+83LO1Q5AwOIvBloaG0ALsAJJHRM7HR6yrCOk2zQwqdPTmSjqiG82Sp/3VawA
Jx3hvhYr/2ekRL5H+SN6vzX1xHj/QQrikXmRh8Hs15z6GrZb2+EuZYYL32vAQE6Z7a220GYpAj0W
vzBu6/+sS/30vpru2HyNXL3RKPxJ1ipaxQoxUj9R0takD1HxmLtAjBbsvsvQWsmlsCji8YI81PG6
v2o1pZaRfrnMsTZPNFvXOfCttYQAN7AQ0rg2lmbeYcrPQXBfgOy10P+rLtvfYk8pVLuFwJXDGLet
JB0c/wIRMuSsckYC6TJltUgHJAZYketIYxVYDDgMsFAKyS94pGpDUIWQ6mvcYyTn8i9iXY72ca7i
eCkquFKztXI4dhJUOPn53p0XdB3Ahftg8bRu7ysF57R+1/KTNVgYky7zhm2M9/bYJaeHmkTLNVXv
O+90No+O5W9Z/12hotEfiYLqIa2iBLXgr/REHYXC+XAcudD0pCKipmc4EWjt+zwKGpds664EiGee
DghR0nl+MUkN8KosA7FdOzHFHponzrcc/nskT7dO33+tzC9l4h2PYK1DR8IGHcfZws48PcRxvSCt
+uoGQgRlWntEtrfvK9sikUnLClhKRboF78Y0o5ZWuXXBlsf+hYfzDBoKznsQ57ZpOxUau5vGYHkh
MZLphjPRSmQhgGVBbdIt3RrWAKrEcZtp3ewcs7Ydu8FnHS3jbL5jK8NsfzXbF5ptX/BaeVbiSBmZ
++T2KxSfzSe8AGX4S7TajmMb5EFHbqUugiiUHkyWbV5L/NEZQLW7S0qkY1/fG7vyAmHCW60J+Hhl
ZPSMzTjLnPEezzwaKCDcIM2wHPNjUD/Ohgo7g1dYF+xvb3m6deS4Tur+oBmSClukvd+HfBWKvp+p
ZYYxUpx+beDiqCrPxBZkK8mFE741o+Xy1iPzIIa8R9zOlcSxoEx8VHiF2AJj3b8TtoSxy8GtCvZd
N9M1j/25pW4JWNOmzpwTBrnDXmqr/VXiAkE0Z0zeYYMCuXQqrgQeB4WixUWT6IPGOe3gL5Nps8+V
Y/jnDFmEfArxC2G55GvFA4f7ew8NP01y2fBcFcRuv8b9KG1bkskhvgglhT89gfgWaarFpTiJR8xj
Tx8OMqgR4QjHHeqjZ2a+n+bznYzlhlAfUCMVyJ90zbEL7mvmO6NJyfNZfrivB3kIh9J9R4D9cEJN
1W29sE8d6qOILDyquaDAxDipA0OWwsr5YdRFbPfUBpWpeIyfoaX6SfgRfUWZhg3iTSNWu3p5Cfr/
cCt8bzYu5FxbfO5bWGU8eiekltNP2NS1JPMyrSTXBm6xxcmqGwl7IHNtjPSXSglY/afFqsOspe3T
cFZ+ES6Z5rpT3BgjifXFDig8ug81b3SU2PAPN9Pg8ZrZRiG/rtF8NXcJmA9Ou4X/r10+YA0yEE8l
CdTnQ10eKBu7EI/2EFwMzWK1aqdl6ilN2xzS1cml8dFr3iqBnAknZVfkj+dgeMZBSzVmwC4hismn
ILMDR9ECZbczLRNvJDrqODSjCIA22snKmVdoakLCCH2bGhCt3LoUV41bUIe7aeFrPZHgjmDclchI
JBUbIcNOpK3rkgoL8BzVvkyM+WyR5Wr3eWweklq3TLEhxL+gs9HwSDgWNktgOL38MRF9v0zMOhQO
pP1LsdBuDteEwAIdNGPYWlm+g6yU2oElNz+h/oxUJbUJF1hadYJCsliUMG9xv4fNqOLTxwlbhD6B
qNbHFVUAr+hyysaML+GHBeNCao5N0WQuiPWmEr2EQtbNbmWmXmG8oIsLIeBekNCzrX+O9GW3x2bu
BIPNWVvXxuPSphOeXIpksGJ+TrwvRNNI0172ETQGlZCfkRltX7pYELkKqwFMUaXTlLBPzO4As+vG
u7XwtRNEhvL0EtMzJH+Jx9bJGrYQRcb/NuCcE8cDs8ed8bNePAOH0/VFiaNZscn72w9qpWYlZWFi
wK1LPOrx3NsK7BlhbVjU2r+HZDizRrZXAa6Pt4Kr4jcY9wgKGAF7xrpum4U54VffCCUkJ/S+PgmG
uUvXwDug0rJ/fdb6QJ7F7N0XiGH74Nmz54YISI5jZ2QFCmRR81eTqxC1jUZQfus/5/raj2Fjp2eC
ucOm9DYNuHXITWGda+CUw80ZvIyrQHPtqEHmdUWnwOL+Nqf0ZRriM9Jgi2oIDsEKwKLh66O8dnMa
TDXVBe9ehdUp/UzpkwJ9w1+XVil/3cVMER1IOx7aTpLSP2DqOoyh9ruefEdQs8YGQ9AfcKfo3pab
35SU/f4jEwNiEjGZhBZTSYKkCRT99pwAZwi4Hg66bgnfaAn2bm9ENKXNFIpSlKXIRITUEQwoJY4n
5EZ/GnRzI1xBsmczIbgK4hetGp3ZVwHkBqhVyZF2HQAoMhGOlqNOC0hsSFkXjeImkdItN10lPEKU
GyXsDtRGyHzvl4Tbt1cDt92CYQKsMtU0ns7a/C9yruWhF8TYRlGWdMMCWBaQPf8SZ6nO5sz9IQHI
hsq7K2AoS8pe5XocDLeR3ZZP0FmQCvEiExErezJ7O+Xn2+5xU3DbVfRfHVvVmdOUvw1BZR762o33
h/brci+jrsTW7tT+YhxYmx1DtYo3JcjpH+BGg3J8AeMpzjgd+ncQbO0bzNS8FEusHMTxawAl/5MF
MMy8O5RD+FlNxSSQYUDoPbhQM2+q/p6lX6WekFRhiBtsy2taE87DPaUPZpk0DSPTMiMRjBCHUQMe
tjygwD2uXiOnQ2oX0O6n5NP4Muh8Kue4YYJESswTWs/V0qEAEHIix5+fhtR/0A3LYTpZTwd/YNvb
dofNorv8c4X+S9Cl8bRP1B4qjNYMW6TLvwqhM5B02p1D2Od9z342mQBb8ZpXhSNpUouOrqu20mbN
5PUUVyZ60NrSWyG7sMkH8/hS+t13WXYIx21bkRktRVs7NlBZlA6IgxHofdrMAEzgup+aUlzhm2C/
rAr3iqLqQuizdJtIwZgUstVjEwfjJwCJRq3qvEJfW6sD8KNJa8hxriBc519rl0NGGFsB/2nSB6Ba
zpAiMza61jg3N2JgUIUbxbC9q+vaegLY0cWzen5hgkRjeTRv/lD9poiptxYYTqYUglZ0eX5zYOaL
LP7Xnlclu7OlhCMtM3T30VVmyw2sg6AdjqfliJ89PO0JR3TmhLs/wEtffuuH8Pzzo/c9xbse+rWM
8jYm77UnG+OT9dDYZo9vCBzxhLuOVftN+EWLqT9g/v4FVdyef9ZEI5KjZiS70SiuFj+q1n8hdIW2
iIh1ofW+Riy8BVtvClWtpqczMaxQZhUSCUfhQAc2mFOb1Vav3ISpvT4zchbLgTUILdJwkJxgAEnL
NjJeAL/5FxJo0rU0VaVCJrBjxTI4A31gfeEDIUm5Vet1facYAMtMkChfE4zZ9N8iGYtf9wW+ME65
FTeh8xCMrUZmYbIK+4bixMAeQhocVojE1fm7bWplYxykUsFHFLqKCZtlzRg4zAVd0JbFf2pMyKMS
gtzOgS8nP41/MzwvH+1Nrs24AKkucW/XK5RdEVl1uRWd97Qk1kQxdK8opnedNswLCVDG3wIkpNyv
RdVcx+y1buGv2IZUXbKKgccADpx1zcWFdDwDBv+Br/X3ymthBqp3vfKBgEBhWz4SMWt8Agtvia/w
o61m8c3fwl1MUSbh/xKlX7YX3ACnAgDRhcJ7aVozcGOBo3SD+K57P4nfwR6G+BscV3PXUyJFTcCo
UD12UHtX66HTHW5KyCfLm3tL3GADgbwU8ZVnMwaCcSkG8HN9X3YLLiXRvKFmyyiE+Nd3hvyRjlgC
cXs/b+Yn1eJzpo81G8Uyv8k+aoAwGsGM6dBZff2rQu/49ZMHOOL/PJ0r+cCCMbZlSMpeStaNRton
cSe6cEXeX/tZFY1bcbAV/UuFQQifgBOnLUKQY6D80A6HjeKHt9GwiKOdI+NxRbZmwv14BqeFZKsz
CCNYhV1dRTQ3ADjStxhFwDvi0tzc4CtPLgnLpj7D+HpOJM9XoeU8LDj5cfa/9Klr8kyyho8eUzUR
VVNRR7NcfQNI0H3hDmDAB8qMqlYcQbBD7xZsFE5jdbIEU7cihTDUsYVs30RtrpiWggx5jXhfJ9tE
XpuGnMf7zev40yGSN7FTnw2Uw03D+rh4PlJW2NE5yJ9R6h8fcZbwGol8RRYkDsfM/lNX0RYdlO7m
Mzun1FWeIjKGEnXVGrmlmeu68lZ2fh1IbdKQtbk6Hh4fOObpidIV3wyV1cO4Y2zYpSGNRYLP6K+A
ZIqNGHZepnmCjZ/DoEa+B6BPp9p5qFx1bdJAILc7n5+gxH3YHNw6eKb7aNBJjqO3wi50axinCn56
5RQOnTcsOX8o3+8VHcWRhsNr7DJv5qreoLi6TAJARzMZexmIOBTmHBEKwQuZh+bhve+xEjs0sNTQ
ZisH1q0qVUNYuWKtZojOZTplYUZWIox2DX9hTwKPJaws4FtQhouZPrunZzr2103R8fIXvYD96kHE
U0ruQR1KaoBWUEMlGGc5vlWfhIDAhSOb1MsIOGLM0itH8xadgtqQXUkmjTjdld+9TIiv5lV/B5kX
LygjBPIOuRv+yhHRCvT521/HdXh7YjmkPgRkQIAjpn20BSW0GxYn7UEslSYHl2O7KjaAS7Sf062+
rssnc6JGQbn34K+9H+XsWWxrmLvJgTCoexxHIozq+hp6kdP9R5OUZPb8iRk4/XUqXrjhZ/XwlFuK
zjuWvBEp7Q/+kV0lho2Gu9nNPwL1G5caFvEZs48Qq26xHNbg3Smeg+IhRsFdcv6o9rsd24Cr1ZIZ
Y5R0gPPIfAWHfgAfdzs224oYx/NNKTqqwI5iHudtxe5COd6nli4jIEAeO8ahOP7m4xIB2tXiCeOo
EGWJLe4mhIdvMDsBHWC5zDhpjsTssmsdNJ96xa0q6P15HyRYdgExQiQyj5QkGcKknkXHYCiIL0tf
D+iHUA7TmHho/ccozSnzUeiu/Dwuf1wPkS7TzBPJy85PU2v6p/MdDefYVTJSbNe8flaSreljq5ZH
kye3IaZRjE/GGWbnEZIZlxZxTcRl3yk8rA8aruFoC3SLldqCvLFnHDcmemBi1+8XDzfh5UHL8QPL
ZFmSxskwpKyrs1K8OUjNGa2xRQoNtWOCG+ygUdBaPhlO+lQImlt0XMPa7LVm/zAWf27mMZOw0LwZ
P3iXT7P/iaE7l4Hbttgit9IHc2eNqyby/p7/xP80DBDMtxwq8Evh/YSPV2oxgcYk7bgn+XBzB5RI
Jytt2MS9QycalaFASBqGBFNvD7pHKBcDP/SdP5kV9dozTJ9Ye5sTxfRCZZ0j755nb71uIALGZLPc
QQSyM21DNvCxbeLD6iC78NcfEtZoc1Y5BZrXcnPE7lFP1mzdLJYA9FhpeVy1gRPBc0mRgHwDjpAx
Edw8/CDfYXUm3hkQ6qbFWxreoNCK67YR+rduwDX3swPnltksa/LDwSqr07jxVZZYDECDTgSIXejF
B19lDfY6zpFCvcSHg8LoIOq6DdBSGKrY9OGzknjPnWW6OcxDY+Yh0L66+bEzv7oQjCv5A9k+O6MB
vyxqW6FBe67F/OS2W+bcXmoZWMFip8aJrsBYh6Vcvys/83TWo2+drDdXIBjCeHlYU0EViPKROqsD
FWup2RcSEXz8i64fV+2rzR9Rg9J74AWzx8q8YWs/eZBtyp2ADb0io36+M6v31tIPggNFQt5Ut0yF
l6DienpeUR7zeGU/E78KjbobE23N0maB8b7bOFA2yB/QJNwcSGJ0VUa9wCjACfZAVk8wjz4vJePf
9AxD0YMHYSJ+muSRjkWcIwRoLRBBuVg1KUuIGEx8PStomSiGn/9Nut0nh6+SXoTzVs+8YUcspkL7
bn0wIVT6kV2kNWw12ufbwL9yjakyrohrsJeVyXoZ3QX0vAYsIsMl4TtkLvWxNG+PcPRHwEytSd7C
6NzTSJRXIOIssAC/SItLgUplmtWTK18xZwtckuOFvXK2HPIaxID0ZqVntpvOuzsvDVI1wyJfAmDL
1QMK+QvWAqn6cuw9fyjUmLVhlhCz9QiCN1FAlqovxq8MK34nB4FLzQL5ehYeejOuVkrNZ9oVhl5B
LDOqdUb34afehdXI5AyX9VOn2771w45bCn+wZiN75K5DZQkbeoQDhEbh7k9af2uxb5CjJWyj/5Po
OwXGUXh5hjfcAT1F+ZSmBsdBCwI5WKY5tPPwrFEmzW+ArL8v37oYr1+yTgbSS60/Oq4K0pUPVfA7
H6L8MzP3rrMQ299VEGemGe5LrF9EYTYNdjLGnP7wbnyZkAliZ/eFjOctANgeDzd+mkHEf2F85ni2
375a199dkLEnN/LRQppDtl1CxqnQupDcVWW5yMJ/yOduUAtTvl9C7gFMvqRpxPbLSK6wRiIwKRUN
mb42z29MdhodZQDNeD8OzcPxydO4TIoJMQR1jIniYha9dRCbf04+3US1OEL1S4eH09ESdNR3jgBW
smlAzxiuJ5q7MURJ3idixijYp5SMg8XMIJwQ48biX4gAMo/5SYTPiaZ1H4r7NXnKiW8oKDkHC4QK
GFvGLtx419EovxAOT17eohOQJ1yBDLV2h0Irxpj5ZFsDJHQjJrwG+YFabfU2E3NkYvdbpAV+y+j+
er1S9kqdeSLIDYKCC7cLDZfXxlEPJ6eLc+hq3TxVpHqAWcnfDraeqt3QGB8MCJgZ4RvJBOUV7ODD
WXzIVu3KU9bOUZ7wY3RPiTxUqCJ2Rn2MWzNkB97MrHHpJhk6GluN04NZ8X4C+XUARsm9lae5+bYo
nOLB4Obfq4xiIwP/1Usv20GG4G6CSxNvL+npRw5/5cyU7XiT2IfQ5Oqk/GWrZdW7sw0O348sIckF
X6nMmYRlymzACZUdX2PUqn56w9SpSsHzA0+ivzEMnsXIO+hlyFGHGEjVWpipK1gPm72OmmcuO23w
FzJ4J+gmFXV6cLKOry7wfg5VrUDmvuWHQL1lnK2ous0ruvpTRcW8ZcjeiouwCuZDj+deLTBShARM
jdQ1qKcaRG8FQdkH+MFZsrFQ9M22LoInVQl5LzC+RILad3VZBRrgRk22H8P60KvHcS7NKh3afUii
1qCkrAPYxwpF5n6bfJFTV569JO0b8EX/yp0fm1S3FrMj/6mLxhW4gSzVAi/GKliDyeo8RuNToygK
A2lBCmdhVq/AmvZCve0sNRYn0gYHt5zopc8qsvacstCnqUZ2Aci6b5bEyQDj35Ci6cdhtdrfx7fB
icM4bJdLspLlv28Ks+4Cd0tse5ObU1oF0Wt5rQtSqAoJjNVB7NTURlCfH0OMgEt8+/F0nIFCMMdP
M5l2EUoR3LLwhtte7BO7Yzep4iye0TycdJzSJjWvx/CG1qtpiKV4UfK/ZCGRXcuUEhN6vghBy66N
zulPj9eCUURKS+BfbYs7NAudODD+XW/YZULjEeBkXv8m9aZBa2qfAkEMTvHGHQBJrqs/FeuRPUr3
EkDkMC0qCoKHuKUC1NpPlEi4SSx0TVItIPszMdkVn3ktwwJME0L/fM5cv6wVbb77EKLcA+Y/jhZ1
k377uvnxpbSNAT6Yr7IwAULjUTJZJ/NWPiORVwU6s4gmSo09cRzHlLEBNGgPxoGA50GfE0b3yHtA
LzNxTYnlUB0gYJRAzwhRqlY+hpz6JIyNLDtY1Nfdd+LUirmvI6IbN/9GvZmD58b8qRMMry+A2nRv
lx9Wv9RU1mUHhmSjW/MoRouszA5BIX/l8wY//GN6504Z1ihXxXLBS8GMvIHydVWXPd/np5+nkGY9
CPdSVS2Z8wweXImhC/O9osw/lnCdEqHi7jxVZpUfg6xUHqJ1vFt0cm8AZYP0USrZ8oL8+m/xzArS
KoMY4KGfMDxJ97ke2hFvh9JB5tpj6ReSF4I65FOzg/t8SvjnKxtfMoAfrMlCl23MXHQmLJrR7fBe
rCLLVFtv+OkAevVVxpQ94VyNLqoRvI8ytL0dLfvrCifE2kbwzt+JxaqgZzrzUxIl6r5j5E4tAd0b
+RPDMph0SILfNaewDU7GdMCNbXjZhPRSU8e5ud8ZB+Qne5CgoH2E++AJommim/hlSvDrKUZiEBpW
+IS2ISohXEf0T0NwQB6W6e/9aex82JHpmsViHgt0vgpTSa+lUWsfO2vB/SvcN7cEuYYny8LGVI6d
FAsvZWIPPvfMJ9ifo2Lgggq/gtvE2pu/5ieYMNMFrEgFI5ohN5wltVWoDKzzbtYu9kPkoDMTxvQK
dcRDFIJF7WMNO8lZrkpHvBmQ5E2SWtRshcwQu23l6AdCgmwuhHSHu0zLDjukk2G/lTePWDj5UlzM
mVZt6ypXeag10ys0mzOKoOb2GVU4H/9PsOOJqoTQfTTfQ0RFJLkVXjQleKdVdb2DU+KKz1WbEmNu
EgeZH2vrl4ncPKfBWrdipMVyyzdkJMa2QwEIQvSqjDPsKWKfIRK+/gwFj80GaYsoWfTqX7ZWN6Hn
eiTJeM1Sj/LfX40u988J6dnWM9knaCVX8KVUZXvFXidLM/qKpS8unndiDwezKXvifXEbZ0mLlo0S
lWvCJw7x0x4lzEqGK9tkBJHbWC3lvR2ec7NbUmwF0vHiiD7OMuiCU6fbSIfYgobriX0iB90r9BvM
mLPfwNaDz/FEAx3bprY44zng6WP2x11LxadY8iSjM7Ela1oifR57K9wOXosVK1UjvkxLsiKJogrL
0io03C7XRTGZLA175ZFkT4NO0dKyarx86zXBfFGyJhh2V2VsA6/Vh6ehRJf8lcpr20+JyAjO1Wlr
H+fw8naJ+SEubMuXYnUkZEhiM+9ZY/eyPiQ5ko14mgiYzDI2TsQDxXMsotTxcRHOMMoXI72NHeTf
QrPFg5OtU6KrOLEK/juIopUmHzD/GJxz7b32t0pPz12BViW4cV+upi3TZbgYC+LHKTIsicOUL7bM
d8r3xxwwdmkzycrP8TYwWWL6Wx1dwXkL9LGdb0pOmpGYLeIj4ORuVal/TiGiRVS6KboU0s/4FGMU
yhkPxDgYDeWNiY4MxgE7kRWzPx4/XGx1ty7TWsaL0J0+E5SJQAJyaImWCrIIPc/vAv7NAy72T8Yx
4LveNZivlISGccyh6MBjYWCfFaecfAxSgqRYCl52gBzShTZpgrqbSpBO204Q86ntHfPSVmEhVGsg
30SgnOKh8hmOs9a3bX0LgKqQfe6yf9LIkU/rVPVarpsu53SrafdlbDCEcktPu03VRjEXWYiOT56R
beHH7KYTVaEF1TjjZTNtWRM6EcG1m1oKMuO1UIpzCltL6dZ0LhNke90XW7iqBMvIgaZSpxx2Y6hQ
E+1nnvhLAMr6Y74UkgB9bUGTVuCIEHvEQz3r4U8Hd6XteXarqLLadu5vh/MKDiYb7KIwJBY6VWmu
4v/5Gv699z0MXUDmdrkJrZ3/ALDRgKDxtnmQeoXziJH0ZwzgmB2qTEpWssnW45Nx5XJIl3O9CASU
zuTv5cBWYng5EoHrjgsI86gAl+H28/iky1A/Nhb3TfFFrHiyJvnuD6mT0ZSv6p+LydGogfEhy9Sa
JsiuvF2H4bAXPDpKJpO1+3Fflniasp+D7qSxjI6UF+FVbfR8HjMMYV9UKPDmfRNmojDAwZsWkdbh
oWxWNYO+mMdoRwRgdec9+uSB0LLNEpuZn+HbZVtqg9weKVMXj/zpVn8GqH4e/+B2aEWJTigl2PbY
SUfJTs8ZQKqcCcYaCRd3XAR+g4NMC/0lQ2LRYcFlT8JjTPNZdepVcdDpVxiQ29WBiBEZEYJ3hqEk
YvcThsm68yIlwlIbkASi57xTvsVSmALdXOWQF99XIXy0MI9FcRBkLoqJeB3rCuIEZhl4FAhbCrte
aLN+/CnDlU+iIENZvzcMJTKgm0IXcZQSAHkVJna27NbOZcqT3tZBrjFyS+NgETcG0Zqn3/4UkX5c
r6iz7Dmov8ZjuzQzFMyHzKopWpn9V5U0bSEmScWn5TVuCtC3QYEJrNPF1IwDGcZDmbSHfVy3d20J
zFQIEu2M+We4ZxD4HzDVvCjTQka+Hqzl0Z+iTwzmeGCvli3WheQIemQ2MFCoaLmkXJLSecxnb79t
+7qa/5j+D2C6Zvte4JMw27k7WSo9bMbgk0JaKkw+qnpC8lbpwIPok5bg85MRxKEuPxM6ouC+4437
/8SC6VGUtC1vLFbyb49p8mDQjtwnqZdtFKOG+8tbfRIbVLbYAS981ko1YJeQGbopjcAIPvUTPGAj
7w3uV5D1RayLSYaF+KijT67yRSC9jeAOEqnqTDwXYolZCrAf1V1zL2NO127Dpqwo2WBPNX4mZDkh
aSBz/58oUA8eIVhPR2YUP4qYzUJdar6b82seRfKnNPplrb2Dvar0jsbKu6GCh7/XG/Wh2nPUy5U4
YPlcUt4Haf1qgTqarcKjR3B8z5bx69DlMMlcAtJe7E06G856dLVjLm926nt76iw9Ag/S/OhaGvTJ
tWkA81Om/5XU+Tt2HTsym+EHCCLrbUKrp4oYTjFaeXssIEoHc1JSHS4t9WCAfYFNTOrTNRHUzy+X
a3H/1R2fyIBua4ZJJsrnfbtSlJCiyvdMDtoJYP4tTZjNugYLz61FOw0McjcPmxbe1m6laVplW3B2
hf7Yx2gQxK8bi8pXPBRYIQZogIdudTu5Z5sX/GqU2gAAn3/ws6QuiJ/BwnEF8I1O0CFYhxvhBw7b
N6QO154MweD/5lM2+NdpmY2426CwqVrqoV56wekoBYeLf08Wp7kfhNemjZUVP+DUYTujlIYNcn42
s4rTfs/CaF1jdR6LOGBK/wIUqA9oXAJkPBjnLIgVqLzenRVeLs+TIYbldtEVTUWwB2tKOY0KJiSn
WYPHWb5okI4v6aU5p8Oxpe7RKTGOu5wOxZfmZfZWPJsskd2/WqTcwkFugojWFOmxhJ/XbPBfQJW/
Q6zsBcSwl9XDUqKPx6nLO+Q7KC7pSHty/CWGlECjFvM7QHXwV3wDXNRam/52gkdsOKnD0XhpWj0C
pg43ZtRkota3OFIbhE3p8bbG0xvENv1gGMxoYCAtUTUpC+44kT/gyvmSO7OGNBqSfyBvZWl/b+md
9GZeeRT28jZ3EM1z4czc6qVJk7G84Ao4R4nVqtRysDeRFb1YCkoiVjuAMG+GuItp4eO1Xy5cRcAP
mi5ZdR2Rp6oACpVtF/fvY6oFpxuy+YWmNEAmjYPiNmaOQz7D+VwAlLVXu3uxCevBQ3bGnAtoYIAh
tJRnAtLRXOEHytE1LOgtuoInu3BJU6Anf4YGiI8Vvk5epUCFVgIOpO1x5dewyRDsIIbhcwBh6/0R
Ogdjkh4EgtriYD3PlNeGtFEHf58I9zxqg/RqzL+lJYBK5jIcCkrhCnoNPSujmYeWatuAB/liJ2So
pNLB2Q5ucSsr3RDk/jBH60p2U6Z9ec8oAN6Iio8pzfF3bwZ0IDbsaf2CCV28chDC/2H7+XUKMY2T
UtwV2wGmUd3C9zpZSDDtJOhGDvOOjQiH4avSFNf0kOyDIYliZYQeszFsRi2RnHkzYsmSTEFKB+ly
FIvS3z+UvYG7LAiQ6bzXTBI+9WlW60ZjcyMgQMHjUSCDOeLJucZq1a9xM1+kZDu0OyUPsoWh0ksp
e781AaXPXd+a4cgk/o+7rzmb2/td9lm1nV/K7evlJBvLqmvC/ScNi7/8R24+cn1T2ubpKW3t2bni
7gZ+U/gj/87ynKvCvxZBfpg05ea59bqiY3u9iHX42vgn60q2PMzbqF5O0Kq4F8noYm1iaK3idO89
YI+hindB/dJ2/m+a/WXqpNkSJJoEL+Nc1ihuBJauM4H4MLWBUBBi4gWOEqZ1GAayXGw9RwG5Z9qR
MsC88NOzxGDE7zZpax1VtyBg4Tgr3U5KPVsXSNzuVgg/QCigQpRk/wXwtAE91hEgTcZoXEruSxc2
HJx1M+3OUlb9HFb0nDcyCZdxNUavIYVX7Fk9zGiQ3l1KBI5NzRzhRSsjK9H33iBc4cAwfGK7vGvL
SmEYtYyp8NguT7zlgIYFFiQDyDnWQIKWUlCPRoVDOV1rmtGtcZKOJPeDdbbtAiJFIAvr4fQBnyMx
GQ6I6iZz7205Yio2jZA/4EH7UpU+SOxi9aKVZubnlcqbbbXBUnndqriey5miFKJg1CAT9+qiJxBq
NxInL6cv1Ek4GAoyzUsqPeDr0YqCWn6tPHoHlKap1k81uytEZI8M/ImF7AjkC7TRRnHzsRIaiEy/
6x8H4mQFOto8nX5BvC8/fxrTu13FjQPCqUOPVhw8hwXSlSCDSwP9ia8LNZ2ht/EO7+qoGGEEq6Rw
sdVtjSOlyYUMCwXAK/2Z4tL2Ifkf0Z+nKzpv7rq7rLDnrNg6wWpqI9SuVDUtJ+PzCF8WeaQJI1Uk
Dfwun1i5eJB5hys9VRFUqAvs4Ac4ObYNPj3sL5jLQM4gW2t2D5QICiP3SX0s/ZW2KYmkMYbQXCti
WVVFaV+FP6OhgRqgMeauACJRamrsmcKj94XQDWDj/XgjG0YDNob1UG+PEeTBlSSDdPnCpvQgTlDk
UkSCXtPW1KN45MxxQDPygtwlDqx3yUYWCktbEicgsb4jsNdnUtfLGxPOcKE+azNXnilpuO94hFOr
CMfbF2qxQ0NzcJiANXvl1cswvfzgcGBWrmm5t734Ot7wPOn8Wz5HZJ5TCu4z2ByE7mT8Co9DYmIs
vysCuDi8OL3xtnISCRVuEybivpC7g/1mR1RFqcmzXAFt8BscZ9lZU22KxkD7eLzAc9u2ltT+yNjk
xUeMXW7Y2lzxfs8mM63V5x1q2c42iSxvNlfYnB/XJRUvtGYQrYg6Pf6UOvjLBqEfTWmPmeOvf3fq
5YvXGuOOIRbEwitOjNAogr8fMcz8UL1d6Vs/lM/yibl8Lc0mKFbK2+eJD2qyepQX+V+1cUu1ffDh
7OO9etfmwIFmBfo89KmJd3ZfhObA7J7+3+3IT80TdgRsDi49kz3GmcSGiV8+R8IgACxhqmL8Dcdh
A6+Bp1MZBDeslf40rmboiSF6qT/vUOmC3OB/429wWdBQBC8K72SV7UP5la6lwQCYi0SChfOJMGkP
sLHEoGPDKBWLlNztpGn2l+zZgEC7np2z4FprB6lpnVqlXUvw/7afZH6+Om+AA8TAmAtV/C5xP1ir
XNih/lbeeKdZ9FGlpBW2lrqTgCt7C3eZY5F0qLsyHcA3SfMIXhW4dBejJt70Ns+RZFDryJ1DXGbg
N0kT7DRQXE6Cewvws2+Wz9Ea3+tWt4zTLseyK5I0r/jKayUnCQLZemW04klmTV9EbQyd/OMHVuR3
5AfoCdwNPM+eJBZIYxo69X9TiTrDkOgsUX6Q160dQZb5KEx1vYnf1v8Pe8XXIh2085X00nFGpG2x
JkmP0rkFclc3GPr9B6DyaT/Zi44OMLqqwX8YK7+OreccWIIQsm7SWHl761WsEDTkgoFd4wdC8bZr
0TkDrPmlNI4xPTWOXCMAeh1gmRh5VEHg00GCN8OoUp66ahPzFFyAT1Sv+RFXRR5t6OsXq/PDmWg7
PHUhXF58ZguBPpbxo1N5RB5aoNWek9Jo4JWPjyq+P0Db1ZWrqYJNJD3NyVdJN1+zPSDd1R2MNTqp
MV+kQgOg4ElgIiw4QKe7U40ymsHQ8sPbiVYC/QFhW+kj17MmouSmsyX0uW9Dac2pAmuK+uee2dJ5
XpY0QpzuIHydd586PWtgF5W59X5dSZc0SeuTpM2fIH5TZ/RAzMcso6NMKc/wRCm83RRlKACOA7b3
koyLOUYhfz7YpkGMqSOYY7Tp8illMslLjnBR9RvD8CHX+avWaQAdUKYDOuyiUAzvSsmT4x2GSXA/
sXhT0BRj9/zgL8FLef5YAeXwu8qqjSZtI4x3J7G7ClJCq/e1oOmI37KxHGmP/P/i87RYnZeHKpk+
y1mifm9DtHpn3u+b80mm3UnLTVFkf5qd5j7Cm03dp3D9tO2wciZIGSGo9PNoFEF9Mzx2tMVWCW1N
sOeC3e8uRbUNkbgyU5OE3IsYbR3aVW6YLAH3527o5knE//Z8nJTTzLbTa87spn9ErnE4HaM2KWIX
n/s1U5cTn2a2z4uzc9TFsS6PEkXWRcijMlv+WP+Z6GYuBEZzjj2nu57Fn4F3gaVItzZWgEad/5SP
8jnj/IUec5vnKLV6LqoUohRAw+WpEVG0zjnZLLq5pkUTpd9h7mN7oJ0SRKp18rGttngN7u6Fvf7n
dtuCP7UUESUz3K+Z94mHTlJyr5NTWpt3FtJcYGvKxG+GmrNnNO06pPasciQg8bRxgy/8pLAJ3ORA
SZzzxmVjatXIVi2+YyAQwcYUl55ORf/Bi+T3tjxjKFA0FLMnFiy8d4ga8XxFlNvKHxtppka10+kz
N1WJ8iWtdHAQeFuZd63XbNigq2AVKmXLO/Fh/1b7LXYWazfBBxt49pf583ee4oEtGQIu/9anQQvT
3Zh1V5qdnZH6sO8K0qEe+ExNGVDNKD2RqpQwcHDd6gK4vcFCr051U+CkWrjKw+UMZRBETQ03IBWj
MBfeKik/SLXRGq5XEQMmTpyCVcRKMiwRepnE4DJmWJl+FeSah/6tUNwoe00F/f3w+f6uF1ukOgu0
OL5c0AtQg2ClSzrNKckFYb/ixKxL2EYWg9fjBtWCqJQ+f6hj3ImcEG6ZSFMvkIlNtFzF7cJMFmlH
3L2w+pBRvL5JmkF2X7RSqlQIJ1npj3p8vKJjRXi75D8Nd8bQlXyjKPcFlkNYArUPpZaKLiCEiCBr
80D2gEhWXYDErtIQd35sW6xu3qdenL5+K+wK/Puhwry2O917EMOldfTmA4jA5W2ySOYlkJ8cShNa
7msEswf4QdJlM63iv9Atp7r/XrNE1jdhKP53x5LaNJzfZjpin/GDPe6PY0QwkrAkV340LeOxrUle
Btf3P5cWaxjtD9a4G4Kp/EYh0RIe49fNFQEI7N8c5yXGQ9xQMRdz+gfy3ns49LbthIX+tU7sA2Qp
0VRNCJjAS9QvQigHurkDsXG/8tII9gEf5dYOcbrf412gchadQtX2higYwlcYlVNQWDUvv7HyYMcT
6x//4QUSSDC3icmdoWYlpvpupDJ8/hzjvjMqJZOluMW/KFY119MB+I4rhkztynF+so4ckakvyGT6
K1C67qa+HirZgg+1y6xc/KXnLD/2Y3i3SCTzK47uiQOQY+5i4O6ht3Jv5mHxcedx1BYQ0/+Qme+2
Gg1PYBJaZhkWPKOz1GRLDO4x3qKJ3L4/VCFke1kbO0z06+wqewkRvFlsIwRIByS97jp19o5g7Zue
kG/D7bKmdVE2YGuqpfITpIW1UH6c4cNLyyqjoYAmjRDcmFDw7riIK7RzpprIhz1UgrHFwFB4WF1D
+Nlp0AoB2dDC4t1k8AH6az3bUkeojw8JCtCJrY7C426MH863vtxMRYxqwE6/H6yOiZ/IVtLVMNeo
YW87hwVICorxhVL52vFUdFUdxYJZKuyUAORGIUgb+RBEYuz6neXTOp4FT4Q80vySsHUKC7p9jtaP
BXm6S9PTCSMNbJP1xv0ZvWmIcUlvV/ZLsYjffraFBMpZ7EHKPYIi4KQSuYwIKHQWHj67wwtz1B5P
YT4gmBvJs1CMz5xqI0Ysmsef2oQcEZCkX6Uyvw58xb7QvnGcBhk/E23D322ZLudMB1Fq5BOBderj
HlbyXZDP6ESn2cUt00hkJnOT4FSERYUlncvvnKY+kK0gpHF0v2DgeTWABaigknCMy6xfnklywBAe
k74b8ZFHKyc6y163mC8tapZDWoZyZ3VYl5OcidirU61EbCpdRXErdxnCk118i8+zLLRzik3CiF14
N/KvXyPTMK37RyIJvvn5HNtwJsP+DkLRDpI8b1yFNXHTvvIDirepBQIXLvoftxtcJhw1/cFgsIzs
ovUj0V70mx94RMOezRHsO9qIBYUGhrssIzew1FxRxeWntjFEbCZsIImdJa+si2DEpvHZnbZOOgza
aEcGarr1l4tuCIRZ+fXBYWt8PPa7QDEL6p/td4JUytyKUe3HZh5gXccpHM4cZ1OjRfG+Kl65+Kwu
eH03WG1pLMWjMWmw/YFINkKw1IP3Aetni133m6BWeBnuSKTBABIXy/xkxyTw+GXo2ggXhLo8GvaK
8Wma4JUhzqfJCzys1PmVaSKnok3i8DUZvOa2+EVTOQOpikXx0r+astnpZI0uk5Hxg3QFHS3fEUGJ
3jUGMWKR9zoOD8RS62y/38iuDBB3Z3oCPh+DqblQXyDyWzEr6Xe/4vZu7gRJp36xALGmKT1b1FrA
c4/KUBsVHR/I1Jz5/Cjvo1o1NqedsOR93gmjSw+6mCfh76g37dgZQGbMyMV/zZcSX6YmiOrzQE0x
/l9QuaAQn/23woF/Yh8Z/z1N/l8DbAEVxGGkR6or8wnDCBN6rH0LpRiRWeZBKFBoH69RNlEFC+KL
Xwv4SW5DiZYt/pP8yOsluiKz51v3XPcQU8t0XOA2+m6K+KqjhpJ6z7QpifkXPcA/9n2A0FYrGnFd
nf9ATebQxxKZDfW6IAFhw8HjovQ+rQYW8PVPVLQeCawGeVLOYTBoBHIKLyUp/iSyWJxiYGnmiHxo
tE4GUyRFK8aF9yzW/6BYQrbkfyL64Xa3tsy3RRctnqw8sFhi1B2IqfnamD6U5jIBxhdX3w8aepcI
5s/Kj+Lq4ZURNny9Xslb2ByA2Qo2ZQu72Ck7cK/2iZewVqa4AVsJmC0lFx+6bzoqy7QUh5Dk/jNH
fCp0EAfV4mnSkPobBzVPmb8jczDwofeTgxdM9ZHo++NEl5G/NF/ygdRW2Cl1OMkLYEpLaaDQCf8U
Wh8l1LrLhcGIZfxPK4/FBlLqUazCJMZogPuuVp5o6SXUUeWBfEhmFujB6VMRfyqDnfyqCkQFZlyw
PJXEU65gZfMaewXJbQenS2cU4cnTsVWz9M7ewnubSTxpWfW+G7O1wcbtMGH6pO7ZZme2f6e+4UHB
rQByEDS7wIWIm9uIFX3rQH1uTVaKOUvup1kq6piLi2wbwnppitAQmPjh7iYhHRB3O5+H83AEcVWX
aszvdCHDgqs810SmYEq8iv1bYtqH1rPpN9UfKQZ+afh2q1bDTFOIyZpj5SgYgTaK0pDSCLWVG8Ao
0jwRiwFBFuXv0FcCbiuzfB/GXb6Bi6XvZ5vtJwXvb4gRCCLTWNw4q2NmQYx9A5IgXCHl4y3uO6fB
x1qrMH/he3VD21iqr5fffC/03Huy/30HlHTPXSva2UCH/X89hj5k8+Lr3D3msNBvskKQA7lP353C
eaBV1JcmHqgYLikSlrnO243t6horU9wkiInBHOKLalEVBoBDl4Jrw8LHQ4Mpg8bMTUERfWwXYck+
+KMuFn/M5gtTC/jGLBViUTSJUuRmxTplLnOXzEaTIyjiruENaQmvVI27Q8h5czpYHpB4a1PvzvLN
QqM/1UGYZEHzGnCBUVDz8X3LRBTO0Oe75R/0rtKE1XYQC5Js0b1GqU41aCG08qVIAk+X2TnJR05Y
WtjVFq31Kmm9k5GKcSdOElSfTDBcfd6Qv3OU4kNvmGo+JRCMxrkZKG3v8+G5f1plenGtDB0+yq5H
BTdj4LbSzShoLK9tArxBw3BSNUCpDA+H6Zncq/okfki+Q673E1vIcQ3UVEh1Z6wbriJiuDKJecnd
N3vigHSLPHZjxh4AW3YcOGodU85EfZyhKgUJOpi/91+A+DbBwMSlfxbrlk5lHLBIpc5aS2XEfUaE
xrTjXM0fhyjosTAn5uUaWvx8orgonxZ4HFNQm5KHsOz8c/ONf6cheK1R1n7s9dRla6MJS9pFo+05
n86lUdbC0X/S57VBi1M8A14oQFQNt6QbBaMqUsMLGUwSXa84RIkOQD0Vy2L5kRSso1tFamb59bMV
lCRuzSP89f+WNubJvxaZWA4OZlPWz0qdWRGUTGfnc1o17VmF1DmHGi8vvkRRYN6KcbpFl7v399zv
lNcrtX+dmWIjnA7NRpd0qsLUFDSKfs25LWI/kmA+lnNxSSKa60XmudPoKkhN+z2GdgJcWpKp65Vb
yqFCNgFrz5XrvyW2BjnV/p0iRxyPUhyeSTk+SeItOcrsEkBckuycRa7I5v4UvIojLU4H3bvlDShq
4WoTn/6hUNjJ2f61x56DJje8FCqvTF6EH2ezFT25ah1KXFjlL6IYZzEKAibRGNNGzT37PNGZhaKv
y9NZydqSXrDIccIx8d0AQLQlNC7zbUGrh6iXR142RvyFxWHitNYszTkLcBPcORplJcZTjv1XNrjO
PZumZFEbhFzP8jJ+YPeNo+BsGHE46KahkLnpxLyC/19FwFjKZ15M1u2pwIKrEuCovhCBC+F4jP0R
/22Oc0oSBc27BKNhyiIadMOqLMZiA5hpypgrk6dMOiLkgN6Vb4SjUyyw/V/8skNH/Losyz9HCPtw
FPJyW8uxhYjLq6LkMwpIMTY9G9ubtAmPRL4V037sCHSZyW7vCw13ZKFTZF+1XV42oooeeNP8Ma3u
aqXEoZBwIDzYhQ+zsYoLbee4veBw3t6bIB3NAHuZ8DaTOxz+FEy4H71VZkOmX2YntvjqTZVVQNVv
bLcABpdWujzi/2lKQhds2rHQSPRPskidAVPG/KR9Mn2q3/HZ5EJYS3TtczgRuoGmH+kZU2Q/jEVL
JVFZbLi2/mN5J7atS/3b9cTED3SJ0z/aOk9ij1S0o3gDoJDGiounHhgO/SzJkSNgIgmvLlgwZ+HQ
r+jmr0XEGmwAbTSH72eUUDBFrfvwf6VmqLxQiV46vskrGx/Gb2YMGOmnlxmTG0dhE2JG7VGKyU7l
0IZKvC32KtOXbIzzp/mTEW8PwbhjYVvAfOwR7MRoSuGAOtab6bL9LFmGHyaiRyqeNb/i4LCr+Gph
GY1YoQ216KlHWsgcTDpPCKXJ4VcTLvPj7Wk6KXPwXTgm8mnaX4dgF9b5DnjS6XloW70Owc7jc2TH
nDzJupPpG5AU+wryf9jUC9MO9od/SrI4GJZao5Naz9XoeML4mcVWJmLbuKSoAl/ZUZA3wL4Wb8Qe
AtR0jk1Lt1NsDdq/2QsefJ4Qdqh3mYuIJn1IxnLs0LEP/L+mvKM0kbaEhZgOBf730EyrMUxOEKex
+h5gTD/r9AroomPW4Q2UVs8l/XE9ad0aZnNLBLYCeXxrx8k4HUUMiAa+pFKhc0GK5vLfd9kBNqqD
EUdR/kKHcqjVODdnu55XP7+Xf1IlcHTjCAaiSBuie/ngj7ukyG7hTBmEYo2ZcgrVcU5VoxatFyQL
FYsywbSwx1XT4IqcYGXB7+tyMCnE9YfLr8De4uFPKbfLO/I7P9t8FxyeE3NAF1V1PyeipN4Sa6vR
2yhIBrT5esERaILQXl/zLEpMZOgZZa6iyzrFmPL9CsTjImA/4GPqNuhGcSlYPQxx7vAY5YAJkvzd
ayrlJo1jT/z30PMje9PF171fXpAj/7w4HDTeo+bOrFBhPzqnOvHapMQJ+nONRD7h8R8P3+bkSDHC
3ArRrc3t/RJCNE6h5+BIQ6bTOFruahFJWhT+s3jZeSOjzIWTYGYKRu/0ZbobDfqgXOdDHk5KcFwx
012cdjilxgKqfi17acYFfAPQ0ZklMTHd5YrPbV5qaij1mMTsIAEUQr1u65wsM/4+9eph4xMeR7dn
2eVeTAyfAwVfmpT7YMuS842P2fY0giNZnMSmq5mX/EGNEeox3aFvZxgd6NhZF/YsPDDydVS3RMPT
Egmn82PtAAtnVcxxbW4LhvJ7SDBodYne/yF7LO6xfyesyQvLOtmmY0K4pmK79LYigM3b+eSDlQKe
G5JY+HAYTKCNpM2NTPBGyza6i3sifleFc+r8bF1wxTUJ22QGgl+KIwe19DcEHbEDiO3jMMc7GmyK
rIxmVCvl5r92Ag3yaY4+WWPHm0j6wO7et8VwF/ErRU8OIkgToXueU7kENYISo/YGLYpLk7C8cI7U
UBWzPAo+mJRgUazSGmL+AOx0hZkr8jTi1mnUgoTebj+FMNPDA9C2HtklZAFPqxu37P00+ZQkgEHG
LX1f1qQ9TCXivuKRtBKCEiaXrOJ+nDqZnU/WQWs3aSF2bqcyDlnbuqeNukMqP8zs7UOdK9mlG4mc
dO/gtEagS61jbiMP0rxeM6YNHblkHpxfKKoMXkDln2O6Dx7OkEkDq8rrrNFKZO6Y1K0y1Li/8zdd
Yib0XcRdHniR2y5qrRbr3kWISetQMgQ66SL/dZm+6otGHMNtoqC+lyYnrihjehZsD65HMB2n7vK9
7eOy7yKhBDuwTdpw0WNi1qRkSnDcwpcAUkA9pK/IqJWAvMlZUsxG5vk6kwQvpOIlBZI15DcED1xf
IAho7tI2L4maOkhPq7fdQrbLhQRS/rlHjff33j4dVN1m4C/8xLg5NDBc5tvX0KqH8ysntDVubHAZ
kV1v5ZHsIlgxjDsVa8YB/btX47dhzLa8mxULTNCCVh9x9D60HqqZIZ9otJ9ocxTJLcViEONgqMt6
DowMysQMNYLQD9dV8SqKLuZAKGGyK0UWo3yj3YMj0h/zwRR9UG/uDtOsJ1FiqwRigz1iG8v1hbL8
5r5f6kkwilSmR7KZmtWLcCCy5CgO17B83Rv5CayolgoC8XWLBXLM6jWUJAefC67J25H1dFFpCYBF
9GSE6MLWUkjDm6FpvuGxGvxsy/sk+qY4Yy+xfMr4fxMA1YoW2qTRa0N2D9tF/vQc7K8/bj+o1Tsk
GsXrlCTghuR7B3HYZ2EJmNcikoyS6eOAmZo70+vw5kUArMd4OLVZmXUwnMIh/QMW9tbaJHJrEprx
Eh+vWPej5CrblDr0E8Fjo7YNjPv5KobeRCSKrrHsRH/nQgTn50nqA4/feuMbUNhY0CUTdy59Daah
/E7T0XBxWZIVrsFhdYvxSPPXuubaM7KaG5oJMbafqyZeDe+JnaZ7iu9Uv6QA07ZEB7gcg60RQAuS
U/FLFfF6YViJ1cQMdNGDcZsPIGU4g75m3nnSE4zbWYmQ6tWDujRlQLT4iO1ounUbnRK+YtsjtTmt
i7PdxY5N0/e0Y1jOoHou5aeILO0PNC0b+Q2/CkCuePu7qxZi0KabHWb8YieGeLaZw/rkuDp5mN4r
QlpOa6YerdirrY/QtNX8uOllC7qbnMNZDPwCjyne1rnz63tlWmORFOs4l3j6qyE2ZLPksKQlcWNq
6hucDq+KliYfzfTtXJ6Dtgk62wGBiNTX2r+OvzPTOcjrrGTXPId9Z9UvAlYefFxDu/0BV6XlzwIf
UJtdSMWlxSEikQxiOoEvD138rcOzs1uDGy+u+FyzkHhB3cPaJe02t9LsUwp5uOCNh0flUR5mkDQG
QGYdtW3p6ZTEApoiyQJte6IT5vfkfp/jbxgui9CC1vxn8e26K91j1IEXZS+GQgG9o6LPebIh9osW
Y04ogSiCxiFbGyYJNfVcyOkTHo7ieq/7OJ45Ozyj9O72lcCmdcfnNwp3xTYsv0ioPtkOVUxTCHBM
zvn+P7nj76YH0CWZH8ubTs5z3M9ZrLzj8G6hOeX/JOEeNX0zKnYFdQEqkQt56rQHeSnOT6b1h19d
844NZZ1OtRErfn18+kKvWh82ENiUykoEPViX91ur66ohyrpwlIuSQLOlUacs275Tqew1rkl6qQEj
M+NMumQIFgYrwaWaDk2tviEtue+4ktRVq0SEWRAgT6jbS8iWUAnx5FMAPOYPhFIl8I/V1QcyrnPj
EzR5qpTvFjgSVwYG2RjjdV99L0CZ6PEiQFhKe5msNGGq/SHzbDZjIIdVJshYNtnaPcz0/eLrBi7m
w5J37NvqbInZBjuu8zzIUomwkDA693Sx0JSYYBe3olHIZ+sHVAAV7qQn9zK/WxFFjzWWfAS62Eyf
ObteopkW3iG9Do/qEgzuUyMWS5J9rE/+jOZ30dh1hhn0TTzfmSDb4BSKTYHhiVGs6IsV6euWgk0m
9BEbYQoQMhjNukhlmTzFi1xSUkv5/JnCVaP4ZIvuC5XbaJJ/IGC0mBWbqQdXkGS5b1ZMjjozZZnV
rmPO+uTrn/z7bdMFiMtJXj/iXqakgIGqgRohVoypgsZ5MeKXNCSJcPHEwEK0YlVGcj/TxZtvN3Tz
GdaO+jKOwWUhURgRJp2FgTJNscDX2dGC4825oimjrqH8SL6HAyG4n4WgbcZ5oVFpWUWEZ5I6PX4U
R2YkmWavwf0jQBC8YMC1xyyWKX5efHHJ5kxOgILMOwFqsAxLh2MKUAq1QoAfmx3DpQF24ggHLdQx
gNnkcRCESDXTP90QYs9+/pkiWYgMVBv/R0WjeFBcDV3XV0yTYX8Gf5lJbOJDExgoMxiB0xzOLMrY
/zi7M5uLBNkqfKhNf7qawfz6KSx6f6g8ZMFMrdv+7XQnb0XSvP+BwerGd8fFckvrC6RC/OwTxoP/
Yhu/erms4J6Fu12BzF1jJYfnChLYE6qc0aThhplhegEaqJ3ZwKdqXeJ+5WjrR9c2qvaaYpnqe5WY
pxpIoHf/q5rvR2KjDjYHD6hloiSBFDyZ5IyoazdjClQXtgBQOuQVXsi2/egXQNyB1v7Zss4ikN0n
aSZOir4PO44l14ORojpGK3HlppMwq8ccNebRKjNdBGksKeP0hAL743qwZrL3mAUt0x0sFUQsOhZ2
JGtbqw7f2KEoCBWTLtVXpgue9KEE5ktIo9gVw8UXu6O1Y6tLuaq3r/NL2EpKlOFrb0knKZ1s3TNP
Dive9/zla66kZSxTeobzSik+C8VJfWUZLgR2UZaLao7Rm5XjuayMMFOPnPeheWDA4nejRH02bpPx
BeR2JEQhOXb5stpXmdkVUhbD9A5GbupSCOD+dhPrc5nPQagThlWRBYSOjt97L6TJIc7S/ycub37X
34e1ejw6goWIxDksEjMJH4X+qOY4zd37wWsr05ffN1aOwwGWPmqa9s6HlX/4cMdHl0KIXrc7Ooy3
OBmrMKl5jKRNd/aDAJ1Eteg1xbLicJ8NL3/WIbVvWc+LZtSda9gJudlPLzWlCgXh/nYvzk3RQ/yf
fxTWptW0Afq5ENxPlEgzi4TrW/n5di9EAeUN1+Wju2qjEdF27rVTOTwed2TI2NRwuJnZnzmB1oMl
Eq2Yp/ZPbUU6YojmzG5idDW827pReGZ1Sls/3fjctJ8mc1JwAfJUGawsHso2lvU2EsnNT7W1QHlI
wbHFhpo/k4ZgqufQ73NfaBJWDrAClirFd1Pl0Zsmuy94sllLZrRBdcjvkMRYQTiQfLzRDKS0cNsM
Rd3Ck60Zb8N6dsykux1KZl6Uc4yF8mjnT9qf+LAIoa3vI932TNf0PK34yZ3P8CcFL1iGKnX2WdCB
gAEo+E/8vhZ4ObXJ785XejDnomV+g05zbxaww0eEv3CoHCgM9JzXv1Aru2p2+2Di2BROaEPesrGK
Aky8ddeS0S7HgdTDhhJQEm+gf+FsGy18mvdz18Ff5Qb4TXfJe21vZmXrZV4E32ByxteSUXWvwZ8N
RRyY8O3I1A5HosI/2pKF/MFD1waSiK/BWKE8010/27pFBV7WUsL5DlUGyEj9sFefEmD/hKMwpCBj
00QYLaHqCMPWGSI1dgw6rTJHp7jVCkecZEsezeniNWFiLi9hljVHzVI08mNqAG1h1nyKy6rzDlwJ
Us5QvJeWOidQQFL1dVbq2xchU473clyOr5CPNlKF5sGCCFKDJG4s8ZshzeHBLkfGxlFuW1LjYumo
tio3WoxENSD+4QB2ohnNmSWW/cfTk68JtddVPtHCXhlaP7DETvMz0OfeLWNGI606K1shyzTXMNkt
7v3CPZThY4zuZYifPFNt0Ay5gg30mTscx6MRIgdHdaamZtZaNcf9X8fT5jFWA1JY8H3+VDXY+J6J
5zDnUa08xNQp6IeJEs/IgV4aLRgYrQ7G8wOICnuk3pIYoe7KAJIZMRvSyjmWCRlhUERrqlWXXuTQ
fT+b1IZvEnrKny2s4LL4xe03fzyx1tkSG69MU5SN9RfvqKCIEvGpIhxKIp45gK82eGyb4zKZZBUT
joUjWJkQ6tnM1wVS/fwyAgPfyJMSUAwibYB0hmeSdsXxR5PYiDwtnCephXJ+XL2l29u3W44KBIUt
BX7qg1/voRy6alPpk7ZHgUZ2rv/16epxDQLBCSnMnoB1asxxrMT7QhelHQppdjEwkIuB66A9Fg6H
E7rPMjo9WDFIOvbfL4GjlyqJrEbFGWDHiW2bULLizJXWJKgbuEI5gdtorztwSF5+f07VkV2TBwjo
aOAV6I2LR1y7hsdAfCHPAlEeaBQZzyxiBehXJOASsiyX8uQFwDmE5fmbrJp5xbDSj9ZxlWegR9pC
IEvBYqBYLbR7VGWQ9F7fwUBfPr6S72395PjhX/Vpi9Filpuro60rfyeOkh1WnH+2uS6dhKAweEA5
ZgESNZt0lmVMjO8ie1fyssxQzH3SWakIK/cn02q06852KYrGWlGS9koqVKmdvO8TKQ1GOWveSRCi
SYOPHdH70E1SxH8FrBzVWOpVFwxJI2CeoPwd6gkGJJkY7KjKbdBNd5qtd6Z+sL7wzkIEFUAYnryT
X2Jy8ZmkvBOp7LE22w8Sd3hgopisM8i0ckALlYyjOEhwerTWDoSYlo34HsNqhj8fB/ECxsM4GbQi
Bk1wmVDwv+HbhNYOp0Et/++69qeBYN/YwlL1224J+ZGwxSNDjaB7Cui2Sd2IdU9D19FLTjJU138E
HPO5bPgte9V/egZL7rdd97ikiEjMfArAe0IM3dZGY1NNOThv5TrAsXK27TbRQpPQty+oFyEpKgAT
6PxsI1bOGodcR9kYhrap7miTo5X39FhUgta/9TnxmzUl6T1l5z1qLQqrcvNTj2g324qYbXLfVuiv
eC4TgToMfPK1I0ITX6+QrPEqGCqtDd1J5412F2wgIhjVmmt2480JTjEzuhc/rO6sh6FW+n4A4dCq
7TTJ4WP8JAphYcOPMwXMXWul4osD3K2T/ZjrSX5S/8BlzT/WtD7n9vkKLowCd76texhR6iMQ0IYx
CfscSFL1bUpSC9w6uJhb+s8ruTmO+Hmo7chIaCV/7o8RzQJQCKKGxh8kk0J4HoagO9YpQOuXt18G
6LnuCPEFF0SWLWop/FDvXV+JdRCzNfe2YHmOL9VKUFdAMg6HxyO45rv2cegmwXddsFmZlFX0w2L8
9XksiwETkfuDrMc93XUHNBTfi3oDLEVQuL6nmVe4RLaFU3FfTJM34rNaXokzw6+hLHEXAeUvuW8T
nSQbGU7o5gg2sqKJFQ4ZBH/dmuBfTwJRLmPuREz0zYzvuLAaznxiZXR1rv+ewHbE60v70UZnRJmC
Ktj4B7tBw3AihDelvT7NHx8JkzLqY+rJbTSI2aO8z4Bx7Dmuu2+VznX0En4xPOS5L0DFFuHzey9q
zO1EXAE3JiyK9+E4fUop9G1hctWdOFqfx7Ho2Fh7CD3zfW5w/F+lGiuMp6vWXWKwxFa/gYP5g6RA
9hI0ie8ospyBzD9QxLpR6sQUea5qwfJmW5bfhNnk4ig8P4YDsiTz1452aNng1c6HVaLl+/3NoZKD
I5D7ujBSlpI4jCmEzSH/j7sfA5T2z475pr6RhazcQ+Pd1au9grehBZjK4mYs/FIJEuxpzbHbnwOP
ygPk3Z/JQjRxOiAC8Z2+FIVAFqZRddiGAB5aNEKyWfN5OQUEy7D9C0pTISspAyry7upW+CBgBupN
2Oxd1MmsmDHgnTb+tNTGEKMQ7rpG8anVNFaULs4hkhJl53MMzlVdruPdWchLw1NugPSG7rT1Hlaq
ls1AIovwlmT3QBGDaF7418GuNrHnk0L7LxFirMQgVgaW0C6kV6apJC+dz6SHgRaUFsE1SR/oqZYm
6gGd7cEPqLWXXCLYQ4iFFT8is1kiSQ135AabMPD5uYDCQYufK0S3psxImMAZhYgvld/xJU3HaE2V
ocRDIcLiW1uCgyqdypT+3wfwEmxRtrmiGOHJE+8hA9erJPAH69J4VF+8BPtacBvKShDA3kXeBE+C
F2hpPDTK2eIrlTYksAQisfGMaeo1SHtzTU5akAVe8GMRVWwgLI4mFTJ5qrEYkwFbs3P28Ss2y07k
dcYzJ4TfX2yCRdjC7eWOvFy6SMNZoLV2XqRO9HGadzc2K1RHaha5EiWDqV3CtuMDACyGnAEYb2R2
AF5rfC+azSbx+0R6RC5EZAYCPN854uJXjPZDbVQQFWwIqz7J1/mrTScgQK5qO4PrssFyOtiSE6kv
F+8OT+zEB3nIvAhTPw7cIYwxTWUe0fRjPFrsiHvQctrpmcmoLpXc5HbC8ma+MBunxJc2JkUtWtzz
U/d05mU0zkI0ltJ0PyWsVs9UCfdjzdGocXEc9rmDJnr+SLQ48/cZzupFjQm/DiEbmjQUyvcagniE
4i/aTWf6RaRBCIPgfH6FYHyOsCOtSp5A+TO+C9VBqzKhjDiKKcDjgdRuCgOVoIqwuPXHzeRRVDIy
D++FASXUfTbbR00ot46elGJC2tVIuf+70AYziszzAWU4HRbWrAOW3yYxjI/Rb/3IuZtv3a1z4ICb
essGXJO4OUtXCCmqmArHjsDw5v6ntax4P1K4LXcSKsMiwucR1se6BL2wPzV74Ec0dDWp5ALjQB6P
YZBQWOv0AbHCtCwSkFoTdjkzMv6KxmIiCuRBk9me6mchB/DMmhyMY96TrMGedmSeuPW1HNfWO/qR
tP77Ni8JgGoQ8OFhBO19fVCiqJP0kDYDVkKqA5brTVYGEsJj2jzxGfPwWJ28+sMh8r3IBX4Oy26I
K5J/Z6nTCXSoAPkUE9P1yRXS/b1BJusEi1ZpN/fKpO/EG/O2+gaMFta1TdJ/ncnDyRcv4lQ2iRzq
rM1fAJUvlOBlDFFdwyO3I62md2QSCuV3yjLwVtBAvtaFL6YTphkbu3A3h8Td9K/xsz7byyFXL2BY
hb7VJ3vqwf7qG8eOt9sdYQZ3ovlFyvqGi1Vv3Z9Hgo0hN2gFEAFwlRrSb4RlRrqfmA6DMgen2nkW
i9N5Q/ix6J/0r1LqW60okMV8Vp+ZYekft0XvCvhZbmUl77eu5Wz9DFOooZLwoL3nkDCanpla9TUa
BYOujMvrh5ejRtPyDO9+88nbRFV+V5GC/+XtF54trzTcDUQyAJKNatBQLMVhhcqgo8F7tslrVZ3D
CGdmKeJxh6X09K/+A/ZNvY3fegZ2506O/Ji/N0oe8B4pJEfCT4v2z2wbVvjMHnXfkEGHmzu5RX/B
oMCLyNBWSJxdWwV5rNzqEuTqoFy6D4M6Wgb869nsc5G6aqw9NoiT1aLx6tnmgdnEUq86b4SEsSEo
hs9vg+5IIiSs2/1s1++1bfxiMGn81RSsLajaB87MfXubak2YXFK3lgF04ywC3OBcKH1I/q0JM4Dc
M6zpwdb1axVedTu2XxK4NgSqNlsLV6ikDXTGjwaX1V/C/FAkd1iOtEGOVlPvHdK/XQyAbnooTihR
XbJq+h6WN95bgLNGMInv8ppXqOn4qCBwF8d+Lrivu7c1ARf5g7cUrx3LMlkRnCxdf0yBIIhcu1oI
U8HsRCLgi5f8Xgo1vvLtQiaMulCKYlMG34OmtRT9Xhh8ImEAlfHPsRYRFwnNXA4YK/J4HvuChyAd
g2LfYEIqhQHBrt1A3mTZfCevnSj4kq1JMVIiizm17s9kzjUKhMic2FKed5zxEXqRwg0mQR4rAii3
0TNd+zzH4ImzZCQNeq5rYIB3fHcnLuzw44EFPMlhYzSkjllzpChfUlqUY6c7W6Zq7Vi+6JeZyZsu
5oLyAW0PUGLA5c45d1nRdibHdWkspqZS0FV+wOu7xIWcE9W6izpyxCAlzHlaNgEzDUHuuYGHcye5
R9jdCnscq7aZHP92WoMkKLMi+Es01yl9f3izumLKa4hty/w8vop5FTvF6TOV/C+lvmhrhLaW7W0+
DRKHQfN1YIoVb75Qu5YUj2l+MgurSLBCFY3+0Za65ta+yemJrJvBIim7o4GdlOKZMb3Q3UFbp8bg
5gWAhfaXSj6teHsJVjZfBojyHJf3DMTT2H4H53YKRfR/h6LH9THi51QsAvUCYnFehojuOdxLP/ke
fYdpKDjb5Ir87ioeoT/M6CivCN7O3CCUHIrQVNtp+14C3GsX1UC4UBZSYZQKr0VM11cN4BGQlpkP
UPFJUkAEYhAb8d+jOhs1bBu2P/pHGFqzuXL+plkCq08YHDms1Q4Fv/r1qNXx+sSneMM46OMcSNJE
BATHnHYF66tmJRQE5VJB7m6dWC+cFA3GeKOakAo8d07OsVitsIl+StY7mDBwZtTHwqZ9kqP6cikv
Udwp8i7LkHL0TJicYOIrgc8KARlCzRfHXiQMMlMBKbFez5vgxX2cxiVpAJh/qeHqbq52Nhb37mQO
N1WmXuRIqfCgjlTO6feTkCwvCzeDU5a2uHjHzbL5s88cF2upkZHJPSjXYPJm3i3N8WU6QP53ELOS
vqM5kvM5Y1ZmcCVREwdF6RO1YjRF8Xvlbx1+GzNmVmhczAt6CeMmuX17J64BnXNsotVQ3kf0Rx/v
FkTrn4DBgnLBCEYmM7t0VASvj2MZZP8AuxF52cL3/Cu6Wts4jqb8WeHnzAXLaNqMuskdE8yZdAtD
va8ARjhX+s7MtNmXI0S3w9I6SCnumtGbNAG28DOpa81xtxU+hToOaiqA9+Cr2h6BvUKvJE2PCnrb
QWrkpIFJ9UW06q837twZHjOAmEQG4eDkeB1CBdRAbReE9bdF90v+1bzrZUE67cEwtqJWiPMTbLqk
tG7sMNBDw2rmHnAL1u/BvMmFb8qASdJfe11EBI1Np2vGHKKFbeVoc7irDccC89hZzjNb0t+ek1wX
cx0U6251CNisVH9bTIBUIKqXgRB2I1a8AgL7K7TzprHvn7gpiohhWj3JV9n3W1x1NpJ84gIeiNDS
U/dhwgXHJyYsj0I5IZ9grRJdXb8V3peh9zQzEwL/27g1H3xfSzoDhGFbIurDnkxkLiXY2aY/7tnJ
OTWfs0dF6ziwZAaZARLmUnO0XTCKXKymqu8U6elUI2JvwoHlJk5ay+wxjwl3xvE6X0/wLjdjMeBA
nsnMIi//6zcX0dRMXa9+p87t3RYTlun9BBgMQj5gQxc1mBlM+0mkUDWcRDkAa11qys8QMo3m9z6Q
pxzGSHR+ehIuWJX5dVZsHq+XRDf8kabCzOjQsS6bkDtKWNTcQLrZJtguMFRtsN5H1JGl0oqK/ovz
RyQrOx59eQTk5bHAigS34T0ZWCsAMU4oL29UpcqSlkTviI69b3zGc8VOsG1QedhB/pqxI7N/+Zbg
XCBFypiChhO2ukB+32RWhqUv1P47jA8kMLqvP0LPNVSjdIgECbS2fCbRIzXV5aG++ljpW03ktW4F
RHLedvHsLUK/bhIdEOnG3+HJGmhLhu/vRK3X9s+i0WOC0ZBC1KCKtGoudlj+aLxHKV5D1V30TtM/
ipGP1XQFu43kYQJAmT1rMom844BSZz4qKAfdlbOaMOPTpDHCiCQbHIF112ajTDasYAI/+b9odiwl
fzw7lN2a2dvcBkJ6dynKGJtntC+Ni0/Zczphz6xUQmYAZ3u0GxPfMyCvkHunZjA4lmaM8OnNWksx
XCwt+9mdC4rXtyCLU63nvFKfukxg+wUsMIwRxwiaSxxjwMhnHhR9qCN/oXrFVSLOqU8R78TxpP+Y
6JWFUAWYSkhIjHhKQ3swLAcvDeX2yst3l366+PkRJuxlUbULK15nVonKbNnHVdOdfM23desG2H48
krqx0nVoCY78EZ+3XUkN0r0wu6AUGqv1cS1ra18DBBsDJBz0fjfYWFdPTk8VlfAlrDcvdWW0uzlz
OxO2u5FlnMyYqkSiB2hsv61Ic/8oNhTKwkVDNzLEVu/f+5FyLN8mGnzIzMKryfVEVGayFsaMVBPr
en8+0RZan8u1j7hYf0QP8mQRT+5FfTrGaG7g8dEH/PVJW0xGChBQpcgurwC7U7AulpxNfTSx7DYI
BWZqyqFMgUgq3bi/bn91Q7aj6P+YJVzWCJ3OePSF1PmgImA44ouS9jsW3SZgsXyoJgZkIPlZWOS+
ObMymAm7T2AwJn60ctff/1XgiQ0yF7npiUx5GZjMD+KpOsKLRSMSosmhOqnqfDKTvItEv8QfDi0C
ouFbQ1XxSpMSA7abejvDvBUztleSJQ8y9a64fC+pUMTrCt9ggbLNdrgLgMIWWau7dQr9WxIAaJUD
Ha3k5XveWGMb2KL3lB/iS375J7SSuCHsuIwIRdbyx//Y7FBxEmuiPANZodCTU6P785YQVLGzO5Fx
aKQb2urSobspjObTNiR99Mdp/Wf/qxFRNZ9wvW1Lta4wrEvwkCM2Jhp039OJPAR0R+/LrZL9Gh1X
tMVVJE4hTN9ksbzFSKVH3GMk07cMqzB2HoDUykEqO6gQ8YKV87Q69Bz8va/yFzXk3hVQtmR7HggF
rl0eMQechjvoHYoQQsTRXNsDkTDUXMgpwAGrbUA6GzRAzlJO6VDUWqHCrpt+NyJLtoJNMoPIkbyr
dSKza9ThPYtXulDnJG82ewjUqbEnhvr4hGPX8IqI91VN07lOIOalz0CkyDcFtRJIiqHQ44r3Hrqu
88BBYd0vs1EhA8JGu/fjc6nUg/ynGxhE+caPxrbjvJgLYY97m4WDmb/AV3PAFFk1ZeovygFY7Zxi
PB0B48FUbaLBUubs3ir116sYVmghc5gsE49PGuqPYOLuN1xFNCsdgwAsEXz3oPb6tq1ZZM//NVMI
Zi89yPF9Rb6tNzQFyOvppihSqlaWhvs2aJ5+t/J1Xxb7grmXmGBrOYQE/gL3JRd1rjX9HtR99pc4
BZcEMpQ2tVGpnhzeWAZd2ClbmbovjmlO8etyGxTTWuiAwHPaadCQiboNvyCvvShWcvppgu7gstqw
Sf82lMdAacx+P0xlOJhJRPFeg8GHa2FN34rLYRRRLAsapJ8Kceq4gR05Rs6Wg1qO/XGR0exY5c1k
i09qT6Q5QPJ3XUHeWN5Y0NrLG+SZ2cWbxygFYXa7Zku8OB5bRaBn7DF9lK2BWh3MzsW0VOCedDO0
GwMXhc2wq8XccceqCrio+ej66SlCdZ7GpvUQ2I7wUNgdiPs//Wy5YIxw1hauhJAUCIMPNjrjVbiw
1xEdY9fmwhNJQq3cy+cceix4v2Xa7eLiALi5mYmoyXhDurOMKeQQfHJaojSw6NYSHBB3E/hlJL8q
S3p9O7EaW3E7vu49ucd1lfvTzMENagienrzL37oJdorWasKXJ9PHDQmRjPtVhU2tLVVkxe5bxHt9
2yzkrtQ1U+vHDQTvyciOqIG9hb0r+VXAitiTCYrAfz+IDV9FUh8C9DoCkZZQp1gYrRz3lyw0Vit+
TxUYGhNt6qUdgXTsdlJQlrmRNQaXmOBtPxXQzX0fu0j1GBbUu2+eS9ZevcgOl1gvrsPomQNZvanY
/nTC+3z4vFUmsjq2NFx8zyErddNlh68yZXYL9jwB9nCA0E/izKC+2Il1mn9zoVC6rRVxjxs/Yvb0
cbyzQn4WdzY03Lvlwrhl0F8KxlL0K4V3oYD+BOvb+kUUiAdhLt18xjZpjHFGNGZzoAVIZVDDyji/
ImW+xjfS07foI3KgZy9q7JA75pUEeVe93gIji3PTL8tYh2wZa/vj4TQWAMgRYrpZTnDzMFHEy486
CBiaNiJaChJz+/gK0D0QDU5CIfBEfjEcaYscFLfAqh09K+yzdYXo3ElweEUcShIndf7XMf+oIqxI
PtRmoeWSMdnvrReVAaLm8OAxPwdugFtVByNeNIxk1oZK1f/JZrnEVKtQwD30bJgF5NGDetyqd5jm
Rpaf//fX6czjbGhdTT9YjjOvUsYkAZ3muQ1mbElkf5ECiWUMCm5nCAi8KCIaFiXlLAwvUI363VMc
3J0hXLt4bgblr73eAd2ZTTDJ6UN+5YHx8C1jK1EoMxmCwYUfWzmIUbARVawCbEIH/19E+d7Ckk+P
GHZAfDVT5xjn+rqVc4J/ETOb14uZq1VxZSlyoLb9dA4AJzc1LlWFEydkkn1EW72KYeEZswx46Oci
zA+1L+nCP2iSjAn0oVcXRlxqlSDhDxhH4WpXBwMfSLvW2yRGRXEbtS2J/Ldud+ImZ1Jy6L6DT94T
hpymc9R2R3x0N2pUIQ4Skd37IUTTXKhArdkH9glzI1GFSc5/wksA63eHlDUu9DocbvDbwIpJN+yX
/7HUtXMT+XEzGNTV6dzhAXRAAqWZ6sieeA0jTovsjfhfOqPMwSAJt+4+YZ2n8owHVPvZvtA1lD/w
fYwMVNrYEmgfc170qptybEyEXraZSSsZ5uq+Gcqg2ZbSl/VvMWF921T7kxYWU9/F5vnlVk3OiSqH
Ev0HcYZjZxsYV97yXptYoaL7yeNBawvi2GcfLPK40OogL134Yhp6GHy1Ltuxaht+YxfUdSaIM/wn
QYMErNPZSgE1i/GDoNCTK/BYJlwWeLuVp3LkfneiX4oXYiJU5k3/mFiYvHScqfYP9RRvrVna8rem
n5rdL8o14U87ErSKQZyISrMcAWYjdGkKPO8wU8fhppj1Z9cFdcdljtVLCeYEQkNQJ4g7uagul7ez
DDBc1hnBoba5aE2km86ZdzA/43NtaKeZvvtT9I2CqTWEbJuIOkI/6cBdtpvaDDo/4zKnYahG4iS4
aw0lNNkHLeaLt6gm4c5FKOUpzOoBYtlqhntnUXo9dur6XMw57mQ6E8tE5XU7stze8BhOLlpYzxqj
lQ6dD/5elefhuE05KMsL6PbCbz25bwgOduP2+nAGHnDkuqTmAxQMhR5jOq4wa8u1cEkQhcV2LG7o
jHcKHycTjwF2WdO7NNU31fKZQtYX0qWEhLe5D/oZBKGH2ZRdF51DW1Zzv7tMWR1de3Md2V4D1qgh
GTCSAAf6lvZLLG4CNd9ozmgQJEI0s8GiC7w3BoNHujrgiM1DbJXvAZX4k7dPZaUK2898bKi5OmXS
FGfAKf/1KeOkcGGEenpecw8BX1fhLuzuiZem0uANLle/5vT6/keymq7USvWzODbkUnInEsWsJlRd
xEmL/ChUX2T9qN5Xems9fHbeXz/VYtc+JmBvHI8B850aikEEvbb86or1r3Wd4Lms9YSGaS9VM+d8
vR8Q4IupUtb/2BioVvDj5bI5D1u0JcBZrPzdgwl36MtKbCfPfkEG7o5lWYFKgAsqa7zFe8/dINiK
jh6ImJqhNwOs0B9ij8MRyxMSqRMGq0DAr1/R5mzs+1WwJDdWFOn9KPM9SjZ1J7GWtpNeS+jnykos
0FSwGgTsHHRNvm1TFrewaztrbcCVZmXTAgJ1g9XPiT6yr07sBvS66UqVemnVZTtUQ/LXVakAZU1b
Pw5bthsLFzdF0DmYasIeE4DOeRuLlS70Rzb7yMpuihRE5WcmEWH4Zm+0JWZJXQM219XSiVNcTuym
iknFUSEoT7bpPsqtVnyzDDVTrvvkkGijDLW7ficpHXE8om5cFMwYUk4cJLUDUdOayM23KkgSTP9N
FdYvW7t1UPxxfMasZSKiVX/8OmPGWS7coB1LfkvsWHo+LzHUGQmTFwtDtNG/dUQZZnm37XLdBWOE
2IGFmWdxFpcgt7NYoLZNoqyw5xf3KzcHK+5hadlsSjaAd+w7lYYov1gDT7FtJgsgEzHX0u1+PsSt
+gY2vkG/HA5t4XibeS26r/RZt2lgQkg+/5yC/F7Nf50nKQPhNRxLjwK8WXIBZjL4T1jJ54jEKYEw
zXXGL++HrN7u3P/k2jop3pGSxfFDFx3F/2mGGxlJCcCmep1a5sx8QWwfiR2oONwe0CCHYszXrvJB
2GTaDGwOOqDB3xhRakAuh3XepgzLyRMY4oxNqtglAbttSiZBzBHKYkmu5tCQPlMRiZqELi+ufzZp
vttLE+xFyhYBpEediCFLmwoNRjfin0rCr+HbpI4ZRbq8q40BE6ukx+CzHpoa/1W6y49LZP8puzU6
HqyLjVDZxBPLmEUm450SCeiWaHIOH2MQCaR1XGNKDOFoRYkJpc/mGbkq33mbSMy2Yz/scJ42UE9a
iCUbdU6h/hPIPUKYzOqzvhLDWykuuUQexfCNhXdy19dAn/ZGxHPtUveHhyMmujUab9QYN6Pj9wgi
uGvI9lKitgDxo/VM+Q3KY7oY5HccIvEIvx+s+MGY/nKQVmGqHPWdIc2JMlHxxZxYHzqgzxxLiBSJ
JZfTHAuS833/rH8rVlaTY19m5blGtiWU56yTxdNbTO5QXpANCF1oFcpvXsZGbAdc3g7wz2dab5Sh
S5qd+GhMM6L2HiNlMEsMK2XKetC1YhJtwFZWXEx7xZxra/srGoIUFHoyqXD0KllBvPKnvMGB4jVp
bu+wBOS2r3noQi9rZiQjRfuKhO5kVFTQZb7IFro/jzh73l8feMRkuMt1/r5aOew2fxK/a/go9i2W
N3uycFPa6JtCoLtP/0rem56vjsghpsk1+zI9Bq5NZ72SEPrUdYHxxXiNYz1ZWb67V+Y8jdgUFMvH
yJW7aPhZNPH4YJYT+YShrbLFmKPsIZ/gTLvJsFe/sfTrSxlyTAZHL5GtSCXYTywYnS69yRIKeVv7
H6ag3ncfuAHJjVrZGg04gG6N0W/FaFO4EMr8ODtpcsecVMA7CJFdQvSO1PsgWvP8jIJshZyBge9x
WvoOhpSKk50ONuox3bBLZYItEqppH6qjOtjWRtbsu4j17Lq5ohzfbO3hICcRHUG8Dn92sCMlPHeT
Pmsm6+hTSwYHjzJ/Yj11Q4xAwYNM+ZOUvUH531NpXkB+66gb8mMO/+FO1hlrZo9x0pbYnRLcyYuj
tMf6EDuTnLpqQl5B1FjXb7SHlGh9fq6kShAf117V9BPJi4HeGiqJJE97G7loMl9GAD5u8DGpzQHx
DCTPIn66f9NgxxExgDvn+hk6m51zc2N/6Z2B3w+Tlp2wO61VpW0uZLzUNnIBg07L5/FUeJ/6gcIl
W9cm2TxBIJrOVDVVi1+7pVw7lWN+jkovBKdPvaPz29rhIg/vSB5ByspuraHfk7U4iimshlot9w3q
L7aN4Qgha3IEEtmstP7HjrdhonNF2gEyqbIqP490I9vEqkZsz3+Id/oUD4UFIu0q6HqUaZGRrOmg
MXi9wXmQ3U/x33CLNI9qKJjbVo0CW4Yf1Zlzm5FxghwKO3SRAFbdzpkkBWCcpRn6c/LT918TE38S
/VwDkz1VrGDsom/n3Aj+uljkRQraWrtDCyXQK7IvsJit41O6QzSIPJfvVTtX2+nhdjrRMfjPJ4Cm
kw1DvahhmZp2jeLZ1261t8WwtRZHzFwsSdESsX/+pgsGfawWt4Q/q/VOxwC/w9lcGf2hQMNXKtJ3
DBAhUeNqF6+Cg12sYXTJmuFNxIUG9sgakFWvn1C9io8xFEdIZff22AsoUx2FcHv/+kTuZOjhcHk2
NKy8Bdui7FwEF68kR5kh1K7Nz0eWhn5a6y1a/nCMbs8M28m2NKTqZBIFsMRMrjQWrd7m5ULZft72
Uky269NlK0/39Q0Lg2U4bqrwgYcrdTWPdwM2CEGSF1cvxO28MoIf6gq2rXYa+fPBRoMXNiTneEqJ
QAu9uimPHH4Hl7wBtfjDYm8gnv2vXdgsnMqXXqVkX7YYL44Wses1zS1nnd6Rb0rPlIC07bnjwkwV
bz2wc2gcShdqq4g1Is4skJHKsO1+p7m7KXWT9jPLwBB+rzYG0lLy45ixDZhHwyYo/sauviXLeqr8
4r+b/WzdBMW7VWI4bPyAvnczsCy5TgTHN3N21FkuBsf1O1UYjv2tJJwnRgbArFHP6hx3JfdJ03Si
J+gWhqIXk/QKXaNPnWNWsIWzDErhDk2Yg4dQIcqBrhel0AMb8vMaxlAeDLNHLijYpsp00CiAaVJC
N0tvCowlmdiP7LruaSFcB3w+zwanLOxZYt3aAmrlqosmm4nBdgul9yHpt8MgAk7aFnDqDm69ejf+
pdP3Pop/aAW8PcdEwRNF5V3rBurGHsdcoxssUZTqyLNMq1ZRFhVQyASiY+9TksoyDfP413o1XmwX
+r5lySKMOrfeosKRvpcDSfAdUyUfXE4GlaGq9T/JZ1PR9r0UZySDnV+E/+1px7KUMnkBpEdmaFr5
IP9xXoOnQlFqDQ7WG3gKwTeNX4XOek0lxqukdc3CB9dDWRVnnaDLuvhUza7raEhwCV3hIhq3T2lY
Qa0xm6CepDGDcSSRcKGxBTpscYS8vicXItyVbkfuOisWutlOUDLdhkrFPvupCeKbtsAXWYAIy8Om
D3t69mABpbcO5xnmJBEd7PuqR40sLZyhaSiv+JQvLTUDehjmgEEhiaYBa0USVQcdR6XMjPMF3BSf
PeEor0sDu42HA+xlmVcFOG8JXfnc1bN+8bnzZeG8Xaz3WzYHY6NPXTRSOl832IphqL+pKrerPk/+
qchCUdm8lobcR8GBk6gBQLmcTZcz1K3EAVLHWuNAw499GMOTIYdEGCprpHcNzc84D6p/Td2O2afN
TzWlChsp9uum6XyiqEFp0DCWlwlQJCy/2RZYHGCGdQR9XwcU7c1fftWVNsSOiqkRBZOE7N0P6Bhz
Cs71gDk+PQnnntnMgQCaWQ2p7CDGrds9Aydb0MuW3FlmsZJJC3RgnAR7JQwqlcSVyrX1IZObVgGa
8SdN0jbe2JQi2OQl7iTN6cCA0vRUgk4p65ngU+A5I2zxoTL7FHgNlCPcboPh9O4kEih9Lvw96e7f
AfBF+uO7oiDS3VmdDCuJLFOZyxqRfv5+gZu7b4HMOuP5sCOOyMniDUUZSyCIMJ6XG0nwR9mZF7Nv
iM3t66NxtobLB4XDgBhp4QdNgRY7AjLfBK56fOmKNfr0w+E8CrYhu+V4LoeAeaxnut4yXoeyOHYs
e/3IAnB7vAQXFJbvHs6nNaOkitzXl5XwRJEzWbYYa6dLy042WnFuc6ROgLNjLBcnTvK0syrGtOJO
vwXEqeoAlNHVYITyy3M7mvah2X2fXlFj560FJS9U0nl5272KxpKmL19B038+lFkhQwrcYfMsbJpe
RiXQMlz+RIVzd4R+K0GT7F6NHAfvwinhWkBAQ/gebVKYKdToB/qZ1wp+haSolj82o1Qv+rx9+Isi
tBCQ4gXWLEUf5KIuSj9TARXxXYzeny5Dh69M1A/aqj0QaX6mhokF/wY8+hx8+JMVhRzm0LBidykw
p5mFh+I68nuaWYT4UtPWUvHNLElXU4kbsWiTr4QI+QdD2lJHBuYoyqvJgALbJTJwQJT4CGCNIDIN
IDM27zC6dLlDD5t1yZmy3wlLfzUch6YwC7J+WcvKcjHNoYwPEba0P2iVF2H1IEZHMJLqQ8NHtztq
ghRQvyb9AoYLVBabAWQ3rJU9OSF/DWlNd73ybBz9eyUiPAnEYkDydVogTpk3dD8oUogD/lqPJX7+
5CUIg2EpCm/ELdcQgcL+KQsCC2RNdk7lseQq6qwIIPHfwNWP2Fza8hk+AWA1MmxM3/F7FwkIFnJG
G4+OVsj7HrwJRgBLlXmaVK8+S30FVHnRbs1JHBeRHs1ve4Q8jnLgZho5ClhMidyYdr0iCAWD21xX
iKEJxeYRHY+XlSGVcD9DnX1x9j02+cQWGoxjkjEewPLiEZqFgiD6S/q/NatfDQHSTp+q8V8yBKjR
Ri0s1g+XREHF3Emk9xlWnIU17LIRfJOILwD23WHjNiQ8beZtuHVYF811legKsI66tY7K2N/Ex5Ij
iyX8l/HSWZA2cTtMLmhbhAbHFmsu6n72xhEY4Xq/vINYH5lNmy2aiTE3zUr2GKe/pPu87t4vDx/J
SOZhW2nXdsyQ7vOGIhwxvEBg8JWyH2XxQSAOEXc8QLOznBLKQxkff2Zvp4wsGVB925pKU7azRbcJ
GuLDq9O2BF7SuokhyEAT2bZP4SNhpZKL+7qNa39JH1U0JREld7Q1TQCyOSmTMqL0KJ1iqBJfZ5nW
uAnQIaryXPI9KKjN/zaF7T00mXNqUfHq1b8nIm8I4lEwLZmxABs7phv+MoVal7akrPSxThzJuiEN
zKFy+2WfF93efukMscMrWpwTmIIjGv3YJr/zEKAhDUxvlK0/ZUstxyIuhvVPUY6xbqSmcOLWjSIu
okf87a4zWus6kpGaIw6LR6E8pPcQfchYDzYT+bOupdcfDWV3I2uMJNIjaE+RBCgFTV97nwyyK2yc
lQb0XyeGpn7JwaO51xGER/iwytpuvLHYnWKZil9UwrCUK/WgZbGhfCYPMlYTcG9ZBhpg/8QTKRQ+
LAsrhkW4AlWUdWV/3K6MnXN/RFOjm+MbiQYGjD3P0R+RA3eBt2VaESEPmuzAUVn0ghaxS8GwJFyv
JEb/Rzcfb/nWUbmsFbTga4Ub0ZTMuiU6fyaXwFgyz662V8+bgfxqHOsXMy5qoDvXGUDw/IrXUieZ
t46N34umW11vl10cvrRLjdvFBorRv0KeUGDZoRys4EutPXudTawBg+Rru4/RVQ1ipwRoeNh7yo6f
9GSvy/KnZVK5r5vfIgb4PhXKZexC8gKrqZA5KSQeBTKtJfgY34InpmZ2VbgHCwdHuzAFOJgKwbt7
eobb9rkfHsef6/bWwZBJPL70PO6wXO1JWcEQWoQaMjH44kUNrxG1iyezuTW0WovuEb+TsQXplNrx
6OZrxPRTWdrbz2cpIZkjD0iBZl16SQZVizmHsMm+qfOxFSjGnXP44hD9k/znolkpEzhBIez/qOty
2rIJU31GObuMcZrCGVU/pMD2PqgVYcewkkkybKsTm1lavO91HvdhwzuSe1PXIKmTKxBZgfAX4CP7
zYWlws9O2Itfo9Uw6+OSBj8VKT2ZSdnGdJKIjVoKUddSRbhEv5wefTW/QqVuY/u6PuE0DC39JvBZ
ebMAR++n8eqCmDR+d4WFBdlLWxN3o8MleOR1KgT/k0oUY/qzVPmpfG0HnxxFyWA94sBAsns5swun
uWKbPM908+kC7h6CIRn0IONybfRvFQIFJ1W706mOilJBKrboHEwScE7ZOSkCpSQpbcIBIDaYj0t2
w+tona81C7f4tcZvdZkgXb+93dQk/FM/+MQuqkr8H3psf17nNmHm2cnoqKJD6Q2l5gZHtJTLllPa
RiXT1DTcAAXdnh5yNqwoh74w7gLxsAQKBpPDl6yY8fA5AqyqUhJZyRnNRI8ZVg0vrx46T0UGotd4
JitBSxY1t1oD+wgWMHkOEYVKaIOOZEFVxWthIwLg9QNvyuyywvoI/hjulW2ZiA2e5IWuSgj6YnpJ
GNgUMly3vR9O8bWm1g2L/W5y9rejN2p3u1D6qPOf9bEHR+Ip9yE+Ul1uYGLIkPMZtq1kR+KAzZds
jjxPQ9MNyHRMLGMs+kWDTs+7nRxu4abWfeQ2R9saFj24tYNn5wYSnDAtsWUgV8E1m3nV7S8mwnQp
nS7KEb/j7DL6EnaBKNN80l6B3SvoXwz4jYnbH/D6xym4AWSWxxn8s8J5Ox0lfKA6vj/1hYuWFGMt
vQojC5Bqc/H7zJQ6GonTneUrW3HxT1qZ2vyzNnmfaLueF1UugjqFbczBJLNXMsOxKlavGEJgfXF0
QYCQEc/Qpl5JgdLpOESJBMKO7/jmSM5WHwlQ6kPXZqU2ICt9DG+Iqx997Bp5HGgSJ6V0Y8rjLEZM
7F8PMn8coOwjzHnHnLVQ5w6Q1V4MTpNEj9665Dmy64iUslzWiVCg7iWFzWJQhsrNSlY4gU37mhYQ
zR3EzCUUY52gN/mizV57j//Sph3Y7AAS9UQUtN2lzrVBunzLhC/YokvKMq+GKIMr7VebTbO4H1mU
cpp4K29ut3ecMpBdYA/rCN18F0hjl42azRx7yW4ElLC3cVszxgPp80C7VTix5WGG1TUIsz5leliY
56ejG69MGr/5kTdeAc+xkJYg1s+NS8lMlUC5P0Gd/49uuup8d7f4y5B5Ic34UfRLY1KJOI6PrprD
ggv8OHJ2QPsmGwjHWTAQ8rK7kFpOr2qiUx/qTSNlskmMv3/6RSIb+Ev8Ahp7ryldMTZ7jb9bd/SR
uJ/N7ywQCkYqV8J1thtmvyPMvgO5T8NsvpcDhH58TZWeDog5pjYguerFRAigz4J9saUXAboZIc9w
wZ2HDlNzyUndmRQSFd38qUB+KqEGYzOfrt2RXOn/xtYV44mcPJk0ZyMAooxb6oQG9MkaQORvLei+
wEX+2TB1JvtAqn9/xElXBggtwbPtFrwPpzLLsesG0zf/sDg6x/ARt1A6Hz5WUDJ+eKiMEh96raEF
AYupZbj3XAvM8Z6XvcrzOAnVjzQDATtGBbUgfoYUkTXEMbeVUY76Yf5+BFmD07gB0IyGeRL5rOJW
WDmnufG2bXtfCypaKncFF9/CgqJBti1I2bzcqCpNas/gfGNF3rbWbtaiGB6RH5zFGGGoTtCzeMIj
IKT1rGZYnbJoeWb6nlRGM0s0uc1tg22FkZZS+DPdhRT+fpXPY+ElAAMr7veWhN5Mm274H6P/WXoW
hHZj+CoyvlesbNgnfakRfEiSqk59DdqIDYyGgikzLujGGS21MBnceR7RnTN9IV7JcfSfhArIdndl
ON+kfHrCTIQPfciknOpxRBBe61Cw/82l93LraULirAmxHDAi6bs7l+Q1yLuF51yh4EeRBqacyfWG
Uw3ve1QRlDfYdgOmBrQvQLgME5YJttJAbvehQgG/1Sn1W+w0CsLH5Qgc1OBV8dRetOAVKzBbB8ov
Posx25cIFnXMfsTK1lD8O1fmjK5of5FYI4ElKGSbzFddegxREjI3joCeiTWWysTgusavhCph7Xbq
SlGiceBJRgeUiUjVouZo6UZHZBbv85xKTojrZ+hpgB4BuSzwOy1N6Q4Fv9tCCwquP/4SJpRXWr1o
0h6x8PbOp97FeJ2Otzz28kf8RbYj0mCUYsgarBFnEcaVkjGpJZGTphmHF40XJJNU+D04GmeZ88Zm
ZtjT8QcHR5PDOmD/CbytnT0iL/F/BuCHuagO/Lm7J8oRHS1H/prmuK5Fl2Z+KPM1RFmyUXVrDW1W
q8+HEBm9zytu+XmTDa60ebOKpFQmK840+XV1cymW3CcQJpkozgyySqcdi8+rC9FXziymEipVi6sf
vf2/5ax7o1uTN7dyZl5lXgXLdN5ozVzQcc5uGp2X8KNbRFrP3zKZp4H6Y0n3gReMGuI45csUCJaY
L01vYovR8ZNYM6uKXZP2lHquaI2yGQVOMPsPQzZQX7QdityGu3Z13j79qbuunUIJC2l2Q2dobTS2
IZ19TfVVPeg4q/BhUHNt9Ih3Si7uQxvi/inIFoeQTOw4IiQfL0uUsMu5pjcXl5UW3bt/lefMyT2A
dKD/E3N7rBRks83Cds4SKLEKvN82OYOU2TijZ5kBlt9WXKvnlQtcgBTfvB+NgdSaSahTSbXhP/Hf
pzlwSKhp8GzqWGNa55yFks4JXd6z5JJave2gVpj9mD7O5UzTvhA7ZlpyTbj0i6OCOrr8VYjW+d2I
RE+b0oNqc/V4uzlJuUq1NOL6JTH2mW+aIURPWEhurA5aJn+J6sBvu8LTIbIDzn8Sqf/REnp4JBG9
ALI2ClhGG/naeUEqmnZB1a9kzhoHhSpgNob1EXFOY+ceJ8Bxo4L67MoJRve6iSUK2LZeit5WUUYg
+M+aFHfciFjBF57neGEJSGeK0K6Bgtd5I+74SMb8rw1//xgy7DCwtoS/qalT5Y7MSXD4z6aBjCLi
JjnMYiLlJzUPdIyJKcs0epeGAW99geI0ttYJL929oxhNN3QEj8+jbGLYQ6hINhjhheBZGvdUY2aW
BBPzub00lUUJuBvunAZAl75foevznnygFbSTLgeUbXsiG6ikhnjEbz+EPgKWZ/MZ43QszAayUWGm
QVdmzFb804wsLNan8B+ckjozhLC9kL0A3TLcq/x8L41TjUCs3BGnZ+uSF6sdFC0lThH0ZeCoRsIN
3OoTiNXyiOITsNn2xxS+uIELH0fIrDiCZhoR8NvEkC02QOzG6bRmcl0fefbjHzI1Lcc1mUQLMO3k
UV5TIcm+ZTsCOh5b3CPu/W7quYv3Cm1OybEWtKI25XTxWLCIKoISt1FVhNT8nbiJepD1YgA9RO4/
2ZVAWscABW3abQ0wqlg6oA4RXwfRYI3Emo0jFoECxsnhwMXGRIv6OgZOdMJeQtMTSoi/tvOtxKoJ
SkywGbQwDxX7s6T8yMBBL0Nn4bsQUg0OELeU3Sym21F44IaagZ1mMEIx2jXEkec6uEHMKxEF4FvM
5hfAoMPb6HeZsqWuDCzlv5PCxHIiKw9J44bCQAXHVBNv7Y7iMJOjmUY0fxmSrnkp2htc7aSPwIwf
30okmR96bhRuT5SSlKqmCmO+/aNI1NA/LPDYoutDahBghcQAS1rM3yG76hxi1icaZWgI3Lwm+ge2
TPiaht0vRP4ctGBxQDGhVNxk7S3bZjDty7oNbWEfbJ2mMwmHf6oEW6apDfSmgEUf4Ib/pYaW7n59
BXNYrDJR8XVDcKTWB6+1baOQK57ou3uc/Y3FrkWRZ8YLWT5nMTvEoekWvzbo+ZotPMAYBF0d4E6S
h72xykRdt/PXEFDYsJw+4H4sIN5AEH4fI2F35v/Xw+bvFWKmtt3LLp1c7WcUSkJbLT7iAlYBA9BE
UHudmkEQgXeReE8rYDPl8Dr6z/mC8hMyS6P3kledGqUF9HY/6MyvJbbkSS9PkUllJXz/vhkFINQ0
hIOmhcjbTln2nj6YPPJ8x7l7jcKDqTKehEFfKQM9jeCdJjipSvKYwMsBlhsg54CIXXXMX43bhx4M
gt4hWx3nbyFVWoOz/Fnl69GJW40hw1MCF9A4VzGYPim2K629y2Zr+XuiumU4NsWc0COcQKmEB3tJ
6708Rl8g32Ul/vzpdpNNRjyKLJU4+/02eCTh3gs12FUFV+miUT4ukMsqwNiqKn8p0apK0zhI/veb
FenxgINzHI8s9nR5CkfUzmcFVeQQG16C2j8B8nQ6ZyHYm+FStsQNMEynKgp8AD4qs76Cg1+K7YDR
EP1pgSUFxk+0hwJTCO8rIRsddESrPyuMPCVqVGmzeU4EXBXJB4mXPITJf2FGbMbkCe70Co/coo1w
dAKMyvS3qmIixp1pxUXMqIS4wyDW/Fv2M2Pm7vT5XQ5ngByfKaSGEbnP//ooF05KrwblxqTvJZ2B
PVOQq9U74PgGw87QadXCoOSzF8No95tmtzHqvP7RVNVLNx55euQkmnVpT+Mbg+qXfSENaj9c3Klj
gB2lCwgBQa4uaArT66Q2wuUcUHdAWLr62WUsvlcl50fSojPlvRFQBV/GGeboBOFTme4j/uBpu+R/
AfZ8XjPmm4qYkGCqZ84uIbCMr/8y4Lb+wHsqzd2rYkLAh5RmtAX3B1MCbSKhT08yiL/doy14CHjU
2vYBnAoVjozFZZvFXQ0FJbZGQ/BQpMrn2MWwNsG7AxUso6XQbXd5oqedqTdO4Dl+18x8Fkb9iy/5
Sp9wtciyi6AV4RU72nK43PoyVeDu3ayJ+kyxQOADySZNNbzkhkEAs8v/NQ3cYPQRlPr2Qf3z77Vr
9vz20kEeNZtBVXbISBAEP20J+0/JatRBazrYACY0/oea6pkI0LF+uXmgrWjnxVxPDJl66MhUNj6b
N5XbnGqxMTxnUcfAX0dL98TPuQW3UFw62Rb7lPu0tXFw0lK3I5PSlSKQq+ceFxSChbiSvQecjFQO
5UlFfdWifOYVkz+s49aZHump9ofBo31Rb9Dtb/34bI4LP7xAaTcDG2imLbtAHrECqUUNN4TYmPcB
fZrksyRlA2p82/HYWWLDp45wvB4pB3EXx4f3Vr5y5B/FDvaUMqFnI96tpm8yi97HkfV0TLvTbsDS
3px0SjbuoVV0izVDjRPq69mizNNaaTfSBKYzmlWLvKYrIXCzoUVQ+g7LX//Y+vMvE90DqUUtYReM
8k94vXl5wpY18OT20MAfWQg9OXkjizD0oA8nJb5BqeAuRDDNKm+4MuBT83YVLrro5fPManpH0yBb
jjAl8EvUUrpQnsP8GhsUeEL4eIDwcVavWZKAPLIB0mCZXy2xhsEP+83PiW38PszY6+NHTXK+grm7
w6sNxqG2VGw6m8ABMzXVlTp963m6FaJbODVgXaNbO1KGnoFiXT4wB1qSjPRxRqAXBx6ZRsYiyJlM
t5YLEv1P4vuj3/ECJgnew7bMYxcIszhG6PJMs5Q1FU0H8158FRDo4L6FYT1fCKejuYdu8xhI60MM
+SsYTOqUWD+T0nDIEoGPSCsK0i+U9q7SlWrGUIuRMzLU+TjSOI8PygP2XD93efAKvw+mMt+9XpJg
H2sutUnbZJCEV7AkROQnxg4LjHl1N70UoWm23hDu7y2+DCnI9INu1Ao4BDCoXzs2ssaJovfHuma0
h4sZxbyVtEwita0QCKWW/9tU7uees9GUqtW7PEHz//+7UlblCSk+UocKcn7xnyoH+xpCfGTY4gkA
aRarWeWhgkg4BPyF/xRiRZIXlXk768fJPnXvFabYk/X+mEHWuCzGbqyTlcxbChhJgvYEHBtvZlt0
H0JsopPQ2bLei4OHrbjb/4vVmxMgvvMcI+uMNPAnzCMK4L8c4sxcDioi5ShwDw/beIJXiAS8yOtS
yxv5xM5Dv1gXUNsaWn7enHn6KpWzi44ftY8V0mThN6DEY+Ip+xzBqHKEN6VhPrJ8HROXUXlHGEaI
0EzQ5ZkbtLQXEeEofvXlynRVSTVHO6xK1rfxBokmfc3w/zPz7Z3ScL9yCKAdqU3n8XUzyGNptWx+
qnme/4nQgLIsU0CpDrziNsy0KS6lb+OcmDM7sxNYNInbBTwywN3pEPlx2vLRdql3nbq0xSevLXJz
/kF8TBrcycO4ENYUah7/EOpd1qi6qauvueAH8pdYc5lLTGEh5FYP9siEWxl1mdiAjuWvQWxWXmdM
pzR9WbTsIydI9IRDWmsadsxZbsMWDu5walc8H/qUR8cYben3AcwLULOF+ftEOtHgEGN4dYLUWraD
Qz8rE4JCDeCJohOLcW2doKI4AtrmKv9iuJFbDEvobfPRMD5AxTeQfK1w/yfkQh86QaiMrufl0lDG
7Z8xelivuolpm+SPOXk4344GsV2qTliXqTsX/sF3XXCSeU9Z1//8X4TF+NIJ/3B4+ghEKDshYkAu
5viiebhmrBgShWda4N3JwWMMZDjAQwqVR7aiwJtxjHrfCNjxBQdezG0lDQRVrXHoyUoj5tmbGaMw
583nvy974uZGKJbwg9ZexnT8h/29CoezrhKamMYOxo643WoM0cNMTbnEiVTAVoA9RKeTZlBm570m
9brQweDOjEUBT69Mb1LdaxZUq4uYfksJXiD2g4KVHmeohNJbQ4FNfoFUpg/QHxEx6l6IwFmyrfEj
PBtUCRmWOJmnNrLok4TsX0Hha/aR9XPEyv+fIDvT9PiR62Toh3iTqfsNIHvMpv6UxFPG4NilFD0h
mKkdRXSA5Kwn/kHhJagENYtVtBlNPAc8nEvvC1hT/YsI/9JzvhgeFWA1sV0hkwsAeiJdhTk/0i+f
aEyabRXrX//ZhLFWmJUKv/XX2FCCEQFJmYTm5zML92QXVWFGU5Lnyg91I0+F2k0cse3+ossSmy1k
hVYVxGhFjawKxWiqEAEkCtUwDwVCBSFfNmZJibBaNxcizzYx2wDOTECcLkev1DbiLC8BT5MhzdnU
7U3VIcjmt6i2jF3HRJPAHl853DEXKVUWK9WqcRJBk/LkYxLkIr9SW5ELJn5CtcRmlzM3Ny/KQAd5
Ics+Qibb2MeHTqE8SCrhhcbPqRDGX1GHk4V9Os5Opv63BvV1ingKikx4jr5QhMaAJRh1KdO6Fs2S
4k0Wv0NbZHkooJhJoL4HRhTxhG7NWWUgiB2LU109314hs4CGOGuCwIjhnzBPFHM6yYElUByUrPGS
+dINaIWzsyAd5fhSGTGa3D9uiEmCGai3xZZrN5mFt+4J91iaSbF1b1AuHErKp/d1rZ+uJRadDi4E
mLteGZV9JmdVGigegZaPMnI4q3+zg6znYrk06c29ZnrppAz4g4uQ1oldhJOChtmbDbZz63ZexPYo
qa2X11u0fUsXaIURsXN1v8NHbhwT0POHH374lkGI0RhNfEVlsP2leTbsS2i0m6KhYLcqmn1QEyzV
QdGQH8NfchnPPTIAQJ1YWVYSrtD0+WXBNnWiUH1CRMk+rqMCgt0UmeTDqV9DnK3VLfWuMj+xE30N
ZKF5rXWXX74DAn9PO0TcqCazwBPrLuLj6md6Avyhlj3kxDYNGs0u1SV8zO8FHramF0UMHAYqqtH8
kIu8grQ3i+DvQ9rdtuSJY6ccJI3rPqEhMw04FcUyB0sCGSmNhKswtWEjmFmLDV8/rv+6G6mLSvP/
OiqhNR+Ur+QJ1LYcKl6oAaG9YyZjyci8Fe+0YR6cbclberaJTOy8k+ozeHA3s117+wxdOgENeqI7
D5TsiMc4jNMEJxpx2VQQOug42z2bB7jFfQLiNPqRR0D2XQ6gMhjrbP64M0mDluHzEfhd/fIJ7e4F
gfTtLvGHGJbQRqiDHsxRZVxtUgwh0jFW6wMpfWsxNOGCgBubvBPYclcpEusN7/ORWWmo3NuOtQNj
llYlXB4GRlD4skg5JNdG9xV9i3H8sR1NNKZHntJIV695tdFGvtLMyFoAU2vNXSITGfqHqQkDRkrt
5DpME8pcGZJ78Y8LaOjaNKgx0dAjei+zQaTIiIKS9KHvZTdrEItQzqwsdx0PAAQwfjEPC4tn4OJw
JMsiWScsPrzizu6KGcien1xSaD1xgajx8pSacr/1NIObQEldRJ/AE4NSmlylVoaGD9M38ditXuhY
mcgRZk8QPWgnXDbFvyygHzA2mF1n8Wmspl3VNmG0VjqkmxTsBMvdHcl6baqtoGcjYGu9S989NTtb
N3PtDEyNH3eZBFT0BYXE3Msa6e67/FXDF9+A+hHrHrpMecRFa+Ul1cTMfMA7Pbp4Fa0Mg9UvVL1u
lr5uPLqsVJ/bz3SK+/c9gxIKkQpCWok63tDjYbT0gBsyrOrcPEQHUQ/iPnUeDQTNf8JOf23BpP54
RBOBizMhDLFiJig7laOp9ZV0KTrggWmKla9f7jJn55Ubeknr85TrhDZ0fRRdp2vcgoLgGciI0j9Q
l1klXSXk2rMcpHz8f7e2NkU/WJryIECapLubZ5Wunh9rxshDzGmuzW+8YNR0o3/9w19IxbjDBS62
SLUnqlMnM1ZnOf4N0hEM0EyL+XH5YbLdeNsJJzb6hNxQkS8Kdi0njO1sJdjYMFnmIj1AM6cT4V4P
Qg5+Pf7d4/LdISRbNVWaYgWHflglHxFcnq7UVWtn1kOG6M44cpBGRGQPK9GUKNKfbrjdh0jZ6AGL
lTkNlgafztiejcpJCAtddpq0SwRhtiKRVPcMUypvxvuJboLvA6VG1af3eAkcUZuPB0CW70Jg7hWS
BxCtxoFsGxBntUWG6uqMsGBxW2WAvXZEyuxbfxgBWFI+YsFSPn14bZzRxE2cWLN7/x59mv4Ma1cp
OTsm1hIwTq8M7pGoeLddW60cI7LQBZ0tC/yKjnNmt5bJqLWrEU7e4O7Xcg8dwrihGSuL5JaeQ6e1
0Cn3Bi2SpAr1Ku3fFWVY8C359gyBnv9qbsP6yuLC0mMF6CFmEmiSVmt9NJDQp+STLqTBHunzQOFW
Vd2YpUvKSBRhfjohh2limEp/iYSHpWzBH6Ihd2A4ZZgJPaQO695A8Fz4OlpM1XEc8kHPz86FVIIJ
Y4wV6oMxIoxLL6UUgMiIE59HLAl0KMnKAUQ83sXYL1GhBhcIypAL0zaW/YcqHF9FYheLhRCzibhr
Gry+pVFzOe5W6GOiFdTAVvhGldfqZ/Jb1UmXbrqkrp0IDyuQ2SdeOBn1zRntgmSxMJR6Qc1rlB+s
B7gZKv1eEKYmoMr0nPvY4sHi3b9nPfXNmT1LhJRjQXUaduTqwiWI6tJi2Kj1vQDGBUMwiUsAZwyW
Pxp3xIdsBNQ6YKFzt0biOXZcXntUEhE4aJgqPYe2OboRHmuB/z92w5yk6WMKiCjO93wOGbwMiwFj
I0Q82HRsJrWiO5z8UpwPKzfMwjkOLK6N/D9o2KTYoUu0WMM6dtQcNd/ZtJ6W/xwIayCMkAv3aNu5
UWi+vr9HeeeMMy4FNBa/F7M7vt5UYB5/xWXN6T5cRZXWKaftjDtCQ+1WMcTl/C688f/uOc2RfIrn
Z6on8mL2M+do+e8DgiwmvHchq/xnN6Hjf8LGUfb2E6gq0mnwtT04CYMKUzrbosVZvLulXySilROw
yqdFpdDI7i4KZ2gBihWxkotvmZXnXuFZ8HiZPY86WgMEbS268iUNiEuDplzEZ+bNm7zzffHa5gR4
2bgpon1SF8AXfmtzHpRM7Zf4XHjLxI6R4a15sM4VqcYt1ZbLDOd+OWxUj2GuCnNNtb95Py3I67V4
OUSmO/rmQTmn4XMwpNqAb2qpZeYzTuDHAbe5x52HftDtxM6vVJpWVM9MZWIPshzczQKP0w78owrV
k0wspmmE/vzVAe6RcjWY+ep6qXZRwV0VtGWrZzzKr14EvJCridnXuRltf7u/bmesW/5jSuuP/VMY
8xAsIakDK1Towv+zIiR+Wr+WuT8Xu26eBfaZypMcf5D3M7kNBVEp/kdqCMQYBgEZxsN68f2qyshW
eGVEfbji/WFYmT60kPWqXR4WiYbXw6I9vcsU8IhPACuRYY/kByVN37lPIxs3f/p+TKmhA6p1jB3l
69En3ywekbkDCbeqTFcLUlKCUKyr8DWTfvLHCD6Kj5Ukz+FKpwRgkDRxEJplKHcsJY2RPoTz82uc
czxrqLuNuwcyvTupGiDssPYL27zLsSX3TZPpzxER4/cwxnX0dDJ3/dyU9mlC2FViuWwq1J22ooUk
wNamypu7MT6ISPv0q6Oxp7UY0Vv5EE2q2/8wq7w83VRIeS6oO80rNKtLkeMxskEnZaXgpHgT0SaC
4gPO+ioMP5obcRSJxmfAhImsHJ2xvwKq1pCH7Q88xofVZpbwsuyq9FIr6kdWr+e2wwQYM+kwST92
OmOSRAD/h3Ho5xpYkVH96dCussCBWeC0aq6nD8kT2JiJ8qZLRjKs+9wUIHM4PZJn5kfkRo9LxdJg
GyT6kUu6W5OYip0jLu41WBd1+K4ICkIAxH9/cIC80WUjcyrLk6UGDy9uI+ik5n0BgGHKN2K/bwjG
UHFmBiNm1WLA1BK38IHW91hADvZliopJ6uk3+f5ODDcGteHuBwoNP02Tk6yFzXVNjeqRl71/eBBs
7TFhbxyvL7O2RHCeWoqc4Hu9bkYb7DfJSBmkVf6cdZM09V1YHBhds8+9A2eMnd9i9prBiV4ol6n/
EpzVSuPHgs8YOWH7GC2IRY7/1rb9y3RTu2+DSHOLokc79nW6XUkxGgDsiGlvFhyLT6Yj+UlmeY8N
/DGIoT5O1vBe6lZtchAScU7oD/WTpR+7dysylH8DnhRmInMwLYQct7W3kEMG9YfMMu6y9fa3cs9r
kmNgbOqI/Xuc7XSh/AiDJuQkYs876ILtUPttyEO37ub51c2laIbzw6ZJYm9jZ/yUokYQeIzgZL5r
KXljibOgHYUoITCHHJGCccAjxKn5x3+lO1uxiEyBmrFOPqoWDXP5nQkTfvPwFVHYgRar6c6PcbuH
O3j5uk08f9kDyj8RChwQVgcsWxnK42xhRG5lE04uaFe1bNf0SqmvzU2Z0Xutg+9HLaDtmiRts3lh
99mvKJKUEpc2qPOnuUpkVtcKvMVd5YopBkK0Kr4vPaWm1vTg52gZiA3hzmF+p5Ry7yw8oXYx7QhY
OjCj0naPbP+W9c9r27rzd6GnbJv05hXOvE2xWcgPQycpU8P1D8QXjQnwv2WBlhayaueuSzrK+jnu
N4sFddLyqx6Bya5jwjtBat/44laApYL1uHiGDuLEgvWxLui0pXorkickeXenPPcT+Tm7TWbS1Iey
T6B9oBa7Fo/C9O8fMN2GEC6Z3mgM3jdAHcm6rxZFuU/sh7Kj4CMs2ZDbb9Xx3i9R6Qx/BGqW9E6G
rKDJNwcniPc1CSRMKIf5UqOeqP5eV5svMTTk4NNMewggQj2oNw803uybkN2FJj65eaCUz+ebXMCX
Vg7xqNAq7yk82GwZ2yuumIdav/N/fPg5DTt+43s8zApij6LwUXbEaLiXl/TSik+aITTAtshu++zF
nqVqWFRGvh2obIgUMaQ+OkDR8YHJvgXEUECOnkJZdSYMIW6Dcq6rM9Nn5AV050PWKXQfo/OFmBV+
prTXvXzANNfgDO4QhQIZUX+awBhGZjGNZGbyGyxeBGChN6obcfZGj5cIAo7gRRum8N0NpsyFW13v
rpuez4mMl8KCe9ZikXovHYyrIUz8qSRCXJHsYFaIhP1J+ZIExO5h2rM5igWwaI/RK+bDSveerv3s
62mlc4j+Cg0Yba7CeoFNYtQnbUNUjkCnPM9jD9iz/kGMmjCEMWAhqGab0DcP21i28cpTpY3OIstW
kyg5lBGFYCRhispYkjovKa66jg6nIXF1v/K0532Bp3S+WmiQfxdCP1/+MJ6Zqtj/Y1M0YAQk9yOT
koLdRzZKqDOK5kDarACKeuj3KzcBN53y7vDtEtep8Q4zQYL5+W6YNVgVdSnhgEhX9DsnbfQr1XwC
yi0vvycN1RpcnRBDaNYlhldhW/UY70uR9fzhUOuJweNFVa7OwKlll4BoQHxJhPUZ82vzmj3ej+CR
vyMnPrYIPgvqzSw6XBq/pqIN7GaxpptdNvyAne8BSkkUCiF5kuYMbMF3PHNEge+6pttbDBRjcLlC
Z6dYuC73fA8mu6wj+cKBXg+I+VHO080jQoVANJXhgSb36F8RnuYDUjoS/jDD7VXjOnfhkWUjg7D7
qqgkGc9MJjd6JTaM+KKouP0w1faojYi33FCM5S5mu8vT+2e1CArAlg9Ca3wetAA1znWxPDLuDU5k
OI1xQnpwasBM09XBKX9iijdD9Z2TI56REAFXAtxQ9NeIqmYjgcfA+lqmiGHQCSO5WuqB25rdDf51
78wkrZSUZVpoRn6jjuM1wGSaa4k+OZ0ClortgBqw+8L7SIk5eAddeAqmS7K4yiJ/RBFxUtDEAz7E
iddc3E7u+Nh+Eoe4ClkLQ3CSkM8wTNDZ7gI1+mRwTC2Mzlx3HXEfNR1zB3Dd2dnU/MuQRaayKHSq
+Y7NPInj9o1QR3B85IeLOM8DOBqAuxQLVk8HdTFOekK4voGAXCvBiC7qMoFXLV/HNibfVwx5Usrz
cJMNepfWclzpd6xWEi7riosiyVmeBWF/m81JkZHsW8hcbnmYoIKPgl33dk1lKF//9wg5gwyBAIMs
V+4udqR+qgnoftPzFP9VyNjQ17LmIBJfMz8x/3X2opbLNjEdp39OHIbUzpMld8Iee0UfIkLK9udF
kxY13xs3aAXl0oZxc5Cmf7k/0GZ97VW3WuHDRx0ZCMuPd4UssC5+S9uhazKxJPpS55NPafr/fgrs
bd8szvToOao/SLP7Oep8OYuo7jl/ckYOqSfyy9flvC4dYjTmrJI+bwUt6KDouq5YenTTuwcDe5sB
NAlQI2S6MQJbQbdyX/14qf9e/cUPhyowL/NY/JwQQDA/gFPa6j04d0I5a/7DQBeEEHOlz7OE/YsY
PXjtC0ml823f21kni54C1IBPgfvkGERrgW+wLFFLR9VQSzyY4Nq8QpIYF6eQdjCfrZeVC00xBDvV
7bt6Qu+4qREdsD171mPn4hCW6zDaRTrAbP6atn6j7KxdJEM4RegcfbqdrlZnApB27GQBdHeURWxP
zuAhux088jjIAEO3hS2qtyIiXyTZoXjXPJHRr04qK5kbHvAATbGb2Wc+IHGCSi7glxlpi3TRqlXz
P6TFTDzK1AEOTSRFcCVHHl/ay/RM6lL6qnO2F8h9Bqvge2dsSduzu0SSdeRqXuuzh/VuDLnX21/3
UBFnfnrLW6AUFazkXJVumq/TptSz8XbiHfXJJJvMu9GeguGtPDf0sixMB1gv5Rx6aeT62hHuxXwZ
TILOe1R3o8ZmW//MMCq1KYb0TLfO72vXeHQ0WOhA0/7paHWY0xkZ+PSeX2BcOPcfuSMECpR05bbo
S7d6JP1yfLg+09WW1RctaYKdGsrSYI6RX4gwku7LzIC4tA+samL+ZYbgNSk957/AnDEQoIW4veuG
U5VvlQpfwNdwXIuvHpXZf8VGYCd/MT7m9+HHQKPp6BnSQse1Cg9YnuYMH69OSsvxFksVUPgAt2Ir
XblTA83ZGUlsOfJZpsO6UTgA7Kuw0frXzeUvzChQG1Lo92bZESGkDiRvQSJW7ZTAbgth/htJRyJg
fL7ox8IJLw6fkoBpfefa7RrurKy5HZ0cRPCv2U4hm2YdCYELAxHtdsaU/FReymTMo45sg3rBaLW6
yVfCPpqwBYYHsTUitBSPFtWd8AwseJBVSE3Sgghc5XF0c8kzwOmWJ9GOCa7/6yYwoPYM3Nc9ymzD
9IvlS912vWVwjp7P91fdqlIKQhWAJrWyucbI+jMhw0+117aodqCs445I4YecNgMhB9K0dc61jJ9a
9U3Yhql+PKN4KLPwT3w0Xp/0kBtfq0wgY47jxHF1wPGKPVtQ8l1BBEofwxHYbAM8B3CdD6lR4CSm
XOokF9qwQz8iVffRRLtUOx18kEDKReqUgvh3ZUexgLmT95oTjgb2CB9Hrq4b8UQDkTB7w7gy+Kd2
WBKhzrcgbel9klA7SBM4Chph5sllxCCyAs0Db9khfN9ZvB5VQQhxvwqIP176xzad0C+03MoSe/ZW
hQhCiabB/juf+M4E6pfV3mdCZbHU6xeM8DynES6Lc0tbuMX0cy9YGdbqdpDod5T3ES/2Lm7PKP4T
67dsGE5gm8n+9U6cL13gTjBEaiknW5bQgZacjpTG0wu/fa+5zG63oJDno5i7xIAT7K8m4kQ193+t
DQyvYeObSjR1ao57VBFxkWdLIGACMbLIGuSJC8UszRokEmeSsZWFotTsPg8yfL5u9oszMF8+dxJ2
8tst0Yl5pG9M2/aXBn8XsYYndjWNwpujgwnureQBb0HWdmSCKW9rana8scUeXOBkTXK4x/7gLxYk
QODQ7WyjgnfCDgKckNu8xFj4ut9pWmnWitrbpPjd/NLrio8nK/g7VbkRLFe7+1RUfyhxpWAPTfbc
CCFJz31+rWTDD/NqzqWNNT70dYiSi/xEXwNqVzj0zVNFrlzkuFRcylVJoRxqlh1npsN2wSte01DX
RvENk9N1zYp58MD2NB1tyth9Jq1W71c1eJC+wQlz2DqKN/l1kb5jEcMYPiS690eJfjo6YQyd3JY9
aQetQW192qCbPWkL8H06Nm4cqKc4hbFajyV/8prxU5ePuMd6YBov3AYRH5mXLBGvRHgC+W9mmok3
4KSc4duA9E22IOhdUke8KRMhttK9lQ/yO8IsyUjOKQZFIki3ZA+VKBduygGcXlh/VH2rRiIWIWUQ
Ex33+gLXk4f16mEqwnzSxfaOiQhf/9r/H9jb36W2CieQuAwYhtjAshemV3tsHpJA4CuJMFWpG1Tv
GnaRF4I99zVxXMIcFm/Aqqg6ZeDJvhrjGaXOEJV4LrzRSSRh9fOsGHnvEF7bDOgy+gYcNDPI8FJ/
OXvh68Ankzw/W1IjbQl9jTsAYolwIHIoNWA6M/XidhIdLNY5fQKtCJh3h4WLrXV7gD14X24EaDtl
pnCt5ueF3gcmjgy+pFb8pXEkZfrMcvXxIbOh/efIv7Px4HxocCunPMEB5Ir6NlG/4LMcY4o4omw5
mAd7pba67epJB54DuZO62zGPgDbphvqQiDJ3cO8armSKsllgSQ57vOsmRUL+YZqAQnwfIhVdt3++
LT681tQNoShqX1sNE8msy3zr3Yb8SRSjCrDlZPWKlhrRkVMCHUqE0McPXaKXw+zYo92sV6ZioajW
FM/c6mA5GaxhMYG2TyHUZqHoZRkWXBOrmiTXKiS+N9VSglEK0tD58NxCXtNSkPiS1Fl79Mf87XxJ
br7sMDaqI/vgHeP9Wiz6DWRb80NjAqlrEx1TEwWZ2IrRmcfUi+MEmcdBAG6IkpAhYiBEEjBxwGLV
O90JkfFW+7z1ERj2gyQQ3Z2r8qHkiwMNKd5MEJJl/deSoov2zftDctPZ0XFFrZUqYJA6hWCQ39YZ
DBQSuCfBIopIvEXbN9KHqp5JyWnL1ufMeOvI9w3ozGIFQKMx0zMmPTGOWaY6wcg2ul6jSPi3/XmO
HxEXRq9VwElyUBGXT7Bddb2V+vUDMZWV/bDOwdYHOrM9KBndDddXoB8aiN3eVtVx6DC6s2glabK+
QM1RTjo8a7iJ0AlBiLZEBUQKU7TpsPdLNL71Wo17oloFOwA2jjgt1qJYXVtdIpWFLITh8ko/p5x+
6N0KsrAY+t4leI1pr90Tmi8FysLdQnu7Sv5zgRP4mf66ZMuTV/N0uX/DZA+CtFKTflmZbRbghi22
d9dIalza9t+63u/6iXr/ayqy8QQSUMKH4hd9R+voZvb34wLGOYKiFhHCtDF3HQXF+zaEj4YY8blF
yZKYkGtNkIoZdvR71HbheILQcd9kwumkn+8oDAJscGFCZYoxICswZ0dAa5Avcu1B8YXqlykZ0sCg
0MK1VbSkwpCZEWNYkSVS2gbVWcRNs8TndiL2IqJQ1rigmaTDAb0DrWFOYgJY8wokmZ8RASqTlUCF
heWP7iYLwwIAoPs3xuug4S5Sc2TzEEuDkafjOqjYFAzcPc14FIcu2G2dfgKYvK5Ik8TWkNtoic2K
mega5aMfZrp7DGMRCmm6n7n4/5HbP8faq95dlHLldScXmNVy7QoDfdpQAZYzqc2FmXsRKu+OSM1t
bdp0FiL4pa+evMbttArh+Wcwleh/IXjomLAPFl03Qc9+vDtKPAobadJR8ThcRwUpY3lY+lVxwVof
yr+9nPNzfNC1JNw4atKrTekMliPndU6b35EnkgQVZHgSpCqhr/lMp2MTPzatLxzf9zd3SWg5QKs7
DY+3BSNY+9Kj10g3C3NGOtpTdL/4FYqrvp5RYlvNlfvnHz3oyW5hWW03x2XJEuC/wcj3GdXh8x59
wDpYDKhC/tZTel3PoCJeHi0zia9l2FAb1X1IzM8P3xaDfjGouZbFZLeldx9dh4cH3Y3eQeok+3dd
LFcDDDgJxdaZkvuSVD7xR+gJtKUoajplTAE4E7WPdvuMxAoWhBqoxw6diDFnIuQsjykAhtljz5sr
Yf3SjmDLI24oEji+DjraWbMNLnbUqfqerCYHhKY5fWy2X7LtsKmKBGiBPLF3vdN3GZgFej4Adjxh
7TkbG+6SEGi8mddN17Gj+DM40jIjv/uW3oo04lDyOXRYVMEHTQU/kcgNiptm6pBNwPXewjctVe1a
EDQnYx3gf7RJ2ZiLYuxpYD9DfPq5WMpFOen930+Jxpzh0MfTvP+gjbp4HpH2ms2nYkudARo15KPd
A/vVFBoJrIFtWazvrEWRtshmY9HIKpVs61SR2iTuD5yxgbucg8FHD0l6hlc98RCWOR727AicZZUd
Nskgx21ywU4cuicddMGZJlXTbxgeTF3yF4xILfag0NMUbapgPe2A120xbFVhrsY9rkF+ztVp7eTk
raEFwbnJozhqnmkSuaa15KR0tmF/63aD7sLV9od6GjLPxy3YaMdKrFbImzr6rYdmWaUPA6JElEQa
qFYt6kLZ74gsa337NVaoWaH/ga0gkxA5kNLfTHJPWqzEC94ECf9dQjhFyZ7kLiIBdVl+WWsptXHK
EJqzwApY55nqKRn9+zU7tR4uw4OIKAqSN6a7h9MH/WFTp0n/NUE4UXXpJslyYnqgwu6ni5VHC3Z7
DVscoO6KUy4soPtod7rfPNn9/5WFiBm5jpXXGhmNuZ2O6wEPuYWoXecvt02kc18a79NkSEnqhkEZ
4sx80wN5UzbvSuj52KxrdrpalvE/euWqarxwfGmbivd8l5ZX10a4HIBOFYi272nylBYGSEtV85Hz
x5R9Qg1xUg16ePn4H9Dp1i/TWwL28Ns31d2g+pWaBq9aaskz0+ufU+DrJT5LyxLYNyaH64Oqacuy
kkPEqDj4WCzyxaI7ufqreVHTg7SGMKq5/B5QMe6RdVubgUOWIHJZNoWls+XxQaJvi7O5H48O+pJ2
smmN2pmKvgT17J5Amz1Gl1Z2OVJjj2Sj5CDHjNwp/iR7ws5L2aMGp3sRaHyzPJssJfNM1qWCIxHZ
onxChXGdbHbhA5tQ05m8ZdwF40RTeHxC8TeOVovg0QHGOdfW65czgnDUJfRGsEJcmngdAGWtgr3V
cd0hMyYEqQFGHC0xZc75zuUN9Paz8IIGNwuU+Ng1v17JgSYgvc6uAmc+tuZnnVRY6CzroeHk9NH8
JBXhZy/PlSqjlTizsiS4rNchDw54WyuQAj+f7Ieu8/FZStiAZh9qGYTUnTGDtZUTlwgHPoUtLp6y
YdksrMaV/KEOjKh2Vaa9yma/gAkm2ZUhKKysvfMwrwNcOebh8255u8502Fhp86mQXU3UEumvwl+u
F3wu2bYltfBD59AsUrblZQfB2PirA8g98vyZtbVC/JRKvESg0bwU++qdyRxUDVn2x8a4B8X12Sdz
RXU1/UBbXcp+6t+GZf+dEJjW0bA9th78j+z9zmVmCmqS+4U2i2+T1MZJYW2DLaI5KG++JAf2HnnT
MsfzKTO+zm7GIsDV5TmD2TOeD8AGZbz3iFHDAva8hPgbvpw3CQaxWcX+BOhq5vWcFEjCix2oPMIh
rh4RBb8XnCYT8ZYyZizfwsPDlqb0bU6h0Fir/Ap5TT+fWJNbBLVHOMAMOH7HjNeUaJka/+KFvi9S
e5izvjuk71i7RwVfZ52VZX8/YcJBF5Tcn06nRyNGWGEd5K4kU1aAxM+MTkF/WfObbJ5cb2N5X2l8
7fjdznZY88QrkqIkqetg1QuWll5y+jrCCd5rQ910Y2awKCi2AMqZJye1YrUoYyfj6XL3iL+3Kk6F
r/Ra8CaHQz+ybWCMLspzi6l6R6mGa2O87zM6eOKKsgMqU45GxNcblsCU3+r/T4KgiqWVKdQTCgnu
l25OzHqpmWvkgoozS55/ZSVtbvV0SdNhtkxFQAtUAkTECdAkm57G99U/Ys1AnYyhIzUlNkJnqk7h
zhzYSJHwSs905vPk3ZExaeQLhnq4I5G0vxmTcEyEQKC+YSUcc/CMig8jSs5tiyRKD806NLb4Jgn/
MQJ5KRW8hiEVU17iiuDWciTUQ4n9xCmOHcvC3Em5OjJ3K/y5xznf0rAKUf1cPAHBIcP+6UVf8xd/
FcnG5cV6nWhLttCRhf1xGhaFdwsTW3fSUOGsiTO1rWrrgH3HRiQZqFhYQIeCGl/M8aguaw+XmuJ4
RjUNWgRAxPqDpNW3EiCACZsYCwy8URlZKbc4jA2YT/WijLwzQSwTHOz88Ra7ScwxbebZ7rUFxflE
BF56k6NeaMvzXVpdFK+ZZMXc9c0LVnKVfb//N12gY6CyYEmPMtTs6GtnL000q0OR8ZN0CT1Of8an
d6t59V5dfszewkAPsiOIq41IadFYq4YTVPSNs0nj+jDRqTkehYPUP0XJeHkcHLKQqZUmE2p1Zmyt
ORZKk7iLcyQMIQxzTDuQm6/VRlnCXTGEiWcm6Btft5IxzuMjch2sZAFjsoF5lmBfl/Hm4prmfyW0
N5fyu1TUPgUXBg3oIVZBY4oKmJSOVs0lqbcQq1HW5aMj52XbrWFdCvRlsqzUrvhZyOXifNBV71WW
hWbAXj8pLItyffgYdTLhqxACZ727emPYde8uR6XxGcMpWoUral2dPQ+UUuZLqq1gmdG5vpTTOQbj
hIof46KFyj+wivsJ4abwgv/caLl8S9Sam8iBC3apQcYkzVLi5YpcWmjV8M7+90iTjXon1wwuydPd
9rBc3awvJnjMd1V1G6AF8GH8llBI3heYGesiFfD58AbjSs2Ze31RPUbHFbgiu6fc+SvqbNQcnrjj
S9UomAByrBLBAvYzP/8nxn1pO2hvJzMQSBkO8UD6hDPwx1kZhAINaoUPtq1WX4rFKMrxRzGIdMso
U8vfnl5lZG1dkJlm699aaRK6w6ZcBAmS29ZelK9XXqD1k5h3JjuZqzSHbtEaQnoSAP4QOSyNA0k6
XM6eaeeKlmfi9sHRqFa0kH6gm9wX43cVgWMGOfrg9GZIJrBaT6U7+8nQywpqjClSqaUbXVXxDoFV
ucdOa6d4avcZZZtlGKc8daJREtbVDPip+QAWjp8Xe+tkDKAa/4PUApf7axBxSoDOySf5r1vYgZGo
8uotmbSQa4fjr1/wQ0n+qQt2btO1Ks0BG/Zt8gv2gKWPEDR26EAlvFROQaM856VkMpJ/70dA8LJ4
DdmBNVSF8l/SwIHbX2cttcNTvneTekBTAoBnoLtEOth4gGMmBwSrcqzHHAaM1Na+OSkihaRVMnk6
mkC9MverFHaW3353hzKgdShsm3aUbS+nP6hEzT6vwB7WkKDalI5lNM77/Pf3ecuHw5+FcoiEJJjJ
+zLk7nyD8ttCFpVgBc/FIZ1vIGSqSMDPbpmjehzBfof52/hBlEFUWywiXFS1NMAiC68hMYf7Vqjq
EgwWiASzr0BseO7bdIPXuvFKgdOIiYbz185TGxJIgIqo+AELJH9BCe02jxJznkBOFeZvcuSwSshh
WhuRubLAOZz2TEX/Vi+8Ox7ZTnyODNwukJho0tjLUWWb7A3odm1PzYZ1HM8A0dL30LI1y5LaaQxc
SUvn0DqHmTpfUqe1DrBc9b09jAzw9vyDW9X3rUFUDwlv9SM4tg2sHtb4WoRkZ3rv9K2J6J26Wp/9
QR7pTQV/3oW6SwoODcecN9A7TbLR1caX5/Ec3CWwdsKz3Vju6vDgr/SZQDRb4nxxM46BiWs44uDi
iiB2rAZMwaNMNiloY/oP45xwumsvJGkRZv1Szv9lD4N6rDhz/iW5GJ8jKliHtsnXiW0xAWIO3k1c
WFpIAC71ZqX2CssT9GoXsaOGEuyiVefSLT4loM+meADH8OoaTCTogJBaMnWlQ+L+3RcZHrpYEk+P
p5JXLA15bnegyxoCOCa3BOE5tGWOQCDYnXoI4sGtdeSG9WBZtwyKV3QB/Mvr9/0XuEI26eYQOii4
MFjqK7mwzEVQXo+26Q+pWOuEyiNap/znqtyE+zcRxRh6YuJ5LRcc+7bzymi87Q7A8TPICwRHFQrt
UO9xO5fV4gbO7PfDPZvSb7XPuPGcU9kQLvToxC44fUGq6ZGEufSIx6nX6jxEU3+n17j0bWYE7lT6
Uf9mngQuEc6LuKZr7aHZAWCOURkndbS1Cdh2idr6odDOvaDK7dmftWIY9eKrx3CZQK6ppaErALq+
VXfA9klK1fNT2qOeCF2S7tu+ZHmhLN/TaiQdiPLUDhsfuajj8YIdDFXEfB3nelAgJXHnAjxyHyUJ
499gqIiLquzT9SElNZs2btQoG+u4Fmw/eUXmdIYLTbrITVfWWUEiCcS2nGhl3FmyA4F123bzsvGi
1q8eP1ScleEaeC7to7A/wMCD5WO0XDfpG5yKfBhh3dK19fZoei8QvQZ/mFeL9B/7MfH0YL0tDd2d
OPzlwruGBgpwXj11XB5TuSv63UwRnc/gkKvX2sWQPrHI6SS6aSM4m3QIqr4D/AY4FSs9qn7G2DJP
2T3Fwb6TSxrZEIwlkGk96w/8sX4hsm2e3JPZPnS8mCce+m9cUAx53ON4IZPfLaBPZPiZIuSRTUnS
hCk9H5IhZaGo8LqOjr7bU+nRt5n/uKit87cb+MlV0nYjO2hUP/Ysa3AEJxY69VnmpRVnkH89smvO
Ch0Z7BWriGkmI1VBc179nCJgbss/NDH2j9uGeRx9rRs+s53PFwQFlCVraYAvW6/0OKZ9XKasroXW
F4liWYCpcsm52/c/SL8NuMBDRNVpUHVVuPMx3xPtV8y/7FWlQdnGqNiKA2MNug8Zc9WLgPidiJMu
ky1scCQD+51ioGPoohRSSLNPr9QOV+cZM6h56HrX8AQh9H1FVv+Bf8J1CJGQsjocSw7Bev2YHpfc
0dwlEhMFWgVhgoPCgwXvJgT9l9FQBhcsEgosAG8AT3gf77yYal/wktfl3Y+bV32oJ5OtrdlnWQg6
hrM/NPauA0eCxqujT78/Q9m+O8xJpZOhgRgg5CvHCM69dmLimX65p36uLPuk7/qOxY9W7mIiNz9S
G4BY7LaYlF516D7NYCuTiBQQUl9elF3qZ9SGX9uY5WNQVNMo2iE7W+XKvf/lBgpGfkAicQtRHvpZ
goZQniZ798ZX7UyH8Erw7kpe2CYTM6BZnje0s4WWytGsqqbV3YtRc0dcjhPaGV3GtKUqnmxgCDYW
m3aBZUZtMWye+yQVwz9XsC4PQWaqXjwNApg63IizOWZ0/my0PhffsLoRGz05ZpbF/AFv5fVCS2PY
BPms4vrAsS0urnapfe+cegc/WKVvSv6Nl5tM/zS/qxek+Ws6CKOUfyUvaLS9rNIN8PHppNKwRbYE
LR8mVw51Uv5MOk86TxrENXC8Zm5BZUrFapMlMM4EOUyrlGzweCl3LQoeCp8SZLTSItjdLEzdQ+jd
QZOHPFVtQFGgIWlJZRi8zUHkELHmze1bsqaEFsvIBduz9zRj+3zMjDUY4fTOTmpE2fnk3n0lTLFR
d+sOxRcp7haDd3W5+aedVwdpSmfG884VE0YCwkVd/LFFXWpUfHivzDmHk9WdPWc6BHVQE66eJ6Eq
t4eJy3ZnKmULrd0+HD7PLSlAmEYCRROeXHxxZlCaOEDV4Jruxrelpd1V/txJUYxZMCKxVrslDlL6
uSdSBCJLJRr8UizvpRsiaDnY/SU2zq5z/PrpJ4ODZlWwEvftbCTbeCgLgOU0Db6YW5HoQZkjumIK
TyIHf9bvAF2iRwgUS5i4RwFHPYbG0ra2a0+kmYydQxFSi/pOmP0KQ2TB7k6qnkaen7kbEQwvZe0M
LWQo+4bZepS3T+3nLbf4rsIlGBh0CsWHX2hawpRP6ZTjTCdKzRBK+QNe1W/Ih1EARqaAPz8KnmbV
xHPl5WAJLe32JKrhLe4Rqx+UYF8Of1sjlaEmp4jUyz71RGto9iBqsNyvK9YnsBtMyzyqPgDLd4mJ
FqUDR1dWL59APilRJ3492oyuoOiF2RW7U2UsEzG5BSqtaXAid2guoHE5M96RvwR2zyXRavx4C26L
tL4wdMsBLOJgGm7GjXVUW1hYcEVM5oaoRg8XxJlRYPqDdpu6uyTZ74HcctJyCTQmDjl8UJwKBxx6
fIENAdsjDIa46/pkja1mxtXhyKRr9paI6Hn8JKw8Ob7Nr5/H924/DVS/1GZVt+sqrLWF9G/GuWVd
9pre0rw1Bw1qLkOs3+i28/2hZMLpEZoKOa30G74cS1ygoXWmVqPUZlQDQHlrNMsNrNFRjMCOnLGj
/RVhnb+HZLYQ9xi9ZRc2GOzerdSSixKutsXwb7SdfDM+GHXHcuKy4Keie6hrACT1vZksQE5zVqjP
6sYhYlrXXYbR3rrimf3gVNallQVlZ14Kncmejco56dNf/88Y3BKNSw4x/MbOxyohkCIEVC8mQDn0
dMmdC404Rxs++gROwQX/FLzypOPKvBXJAXHvO9GBYKAq/18qOP5zVvusPr01AcYJArZpY6xy6XEd
4aYNg+SdSG9lEqC6IosX5ZnELdsm4L4+IGPap+I3tIqFysIEy6YYNy2kv7wZJOoh1adkSqAdmyGw
3/iEADlXqThAkGqwLSK1Hjk6aSR9TNmNnAK1vchfN6U3nbICUfT+FRyeWEE+y5kZeSx+gj1z6IpV
Bx/oNyJq0eBsV1GLrpVddEl6/qG+/QY0hYELMCpNRJtAHnud7hFYH5/QKR58RfNhrCvYcQZi+O77
8kFf+Yw2da8RS43+7gNqd1pmHEGxmtpGx18BWy4CENqT6+wNvCApSQuHn6pwV5N9Vu/goy1+2y/d
ne5ZzI79RfSiBWIZAxNusNOH+RdMz7zWOBBWWIh7cWwhlU1AF4tm2l4Xi9ssPlFzqTUPsvsV/8jV
LwVGqSgFSKTNv8byVhdQ1k8Vu1roOb40DjA5QXAMp1iuQDAH+TGd9eVIFUK4xdu+HDqnxqDCanZo
AjhvP7Zqfug2iZumFxZVyLMsRX8m/xuSrFUQeuYYfT/SYDz8fk2MZqLxlMOYbkIwKtvhFf+hi5Dc
pk+kJDAWKesxOkk4hz8oV0RtsgedOavYDq27EiEhcgq9ezqs4JBRXWqtORVF/xdwx5/zIQUqPsa2
g/mPMWcsVct+O+UHvu4dfhXWIQonDqFnjXOCfX4Tk8jllPcv9qKTxjZ8kvMAfciIf8ok/aA8c4Ro
QdEdG24j/A16Rnepfm/4co9Ujy7gh40ihf6jMZPwoTIqtxrKDcvG626fxmN5sW4xwSRgoUP+zdHY
CEvEjkf0sBnfLXTSakkEctUaIVwF/pqU4BDYuqcDB7HkKgGVx8EFQcdIwBNq2UvgP9CUNkRwMyP4
Ncs2bFdxPAvI18Dx6XGZQLQDfCO/WoSnriPZEpNbqdOedPymWiIBs48r7dOFrXKVZv+Nz1NsY4Zc
+CH4U4Rgjj9lYvaE6snBnDyNwC0CCNoUVN8ogiH1HX7+FxX7VTcLc101XHFvsfnJa9yclICxzIpV
PjLay7XNtKsmq70U33PnOx8YZPz4upIH0XhZGl+MljaicVEg3eNchzZqcNtegIeYObfZkKUKCPzF
yMts8fOUiBwCOWR8ZlhvGzUcqMBYfxu3lArCrLsteYNq5A6rZEKpqzBZGfHukNiowD0GNL7RzLr4
+vM7ZOA7hAvZInQ4Evq8IymS91sT0N0Jb5hAv3ZEKmck1ypWFpAczAc7xmJGGdd42DMBAQT+LJaV
adEXqz3YqhCcDgRIOl9o03q5eG30Fmk7Ym5oQ5QWJGRj2LqfTSyhqNuZsOUxi4NIbpnWxa5hwYBw
hmufprmZbkfk5U9jyiB6n+utuXxhGG2OfrJ6z0ztmIzcH+Snodm7/A8F/EpVQ1IDLLeh6mDq4bWf
5bVBL5WsaVqpc56dx8Su8NORBzLwjGb9SwifajTVOQULB9FbmLazG7Ff7CESKHyTPf+tlUfsjP3+
u9wpoKTtOsZMOw0DRtq6DvXJ3g/RtWI2BQQylO24bpfBShMI1sfwwr1MibOUpNDOlWXhGOcc46HO
WpJOxEUOm15a966To7HCfIac0+MYhq0nVge+adnrQSlj1yOC7Nno4EjRNBTpVxQT9a+B2qphzdJG
XOvYTj/dHgSm1x8SVHp7uQD24ADnZmuUPynfK86WtLkLse/FAnFB5o6FU4n3ybJ00SN8XWHobtkV
3qP8blWzkcn4yfwgA2296MMTd6tpu3FSydIopDy0li26HBF6JH4LuGNNzw/t+q0xhDA9YBmQ1uPc
Xize0+JYj3wA0KO+grbZVEbsmVeXiBCVkbI/LZPTwuPsPODMDugKcLxWQrqtQLEZj+y4zb03u578
QN3n1ta479qJ5/ctOEC/+WSFOlWEgjGiZhPH1E2fpTPiuW0aYL7CCs9XnpPzfL+hGpem150FahX/
5+UZh6Cxtb7RoZForUFUeu5EyPHZsNZF/SNJi95VNy2QEy0Z1yhBlenjKSaphntmQ39A4oyR/o7b
4ZSdO3rf7onpn6xMm3k+iTl6HWRXQXYBuDF7O5pSqF7TVqfrIe713edE3FdsliiEj4dOzUqCcwDr
8wGQ7ryGMinF/GatoNFfF03K9CIrVjaEanXnWEF2vGbHp/tE8+Vk8R1kZ7RCTnpZ3bDVp4QQr+Lc
PdYQlfz7e1brMYcYCROJlpCpN67n4zXhoaIPakMO3Nv5vV1gU+KUN+QtLIQg55pOxTVUJGEb9LI4
IwO9YzRSLS8Cnzg3+LuPe2qiQ1ZxzTdOzvOgy4XGdFqqFgE8nnKf2F8ct8kmb0STeUVrqmfe6615
ndpwWRHGOIBT4hU/8K/Ym39awwQxcGzl4Rt5lkyOF+k221EEwhOrEXOOr5ssE+8p/7hv8maMOQic
vEwFBqjdL3M4yr/0mWGbi9MhXNmM0ENOTuyx3pvqZmtOs4zbw425A+6sY+r6WAeaQJNFy4JSJly2
m6yg9vkb4CgJJr+df9Gw5bYiEu+Qs6urgYYgzhLT+Zl3lUt68pIvP8vRk6JLbymOVdRnmrxC84LR
v6kTw6QV2PufCLb83aI8irjCMJeeHYUhKpxhMYqyuRR5eHOZeSifnaIHx7ZezPA/12ICbGD6Uy+P
L70f7ByzhiYlth4rS1XlUWij2cIUEnUY6uJdzpE8HfL2mfXkANBjyzUyCb7g80aBXFgRH2RPc4Wg
/1+EyCivmsFyJ3kxXCSIs98GiOykf0rABi877r2dvncRyZJuimKECso1wxGlegG9YrFgnk7zjRPe
AUc82rteTngrlL3uRl+BJMdKII2Fl2YSOCsY8bJThSeavLuLtf0HOZuzo5AmomvzrHSIQItn49cC
BXfQopXoVHZ/4VUjIoGGpvd+xIKvpHpDMR1jl5+/al10XVrhHwS0vMYiaviE+3yn8qjPwvyRLjmZ
1Gd22ycD6q5PyCPELyzMhGuKK/RHK7226IHe0V5FHiyLYdTAJ/x55hC+zCu7J+89i7pf/fTYMoXq
csVHR6OoGyVOj/DxkJUTR8zq+3cFqcMZyBvB/U6rBjPtENf4k5XaOVFcwvKObn6mRyQMJeKbwwRm
VrBWlrcHfd2Ffnywj7bLOaxUXK9iOFEVM7OqxcwgaWZ/efmTptffZVNn0WaZgl+KywFbl9h5bEK+
9Opb3hO8kA5AwO2LWP5eqsn5t5k/vGKcCysI1GunJX3TelG/Vi2gNyGE224H4LTyFktxC4ACUU63
rot2kB7G3bFblYaYpwBghtWoMDjHt6Oy+IuwR9c48b05HCfeBVendzAZsH2DGaxcconbo5OmZwnW
9PimyI82DVQnpFIh1UqPQKnN+DjNLBMNG8+D5g0+ck4GJNJOxfhbrEAiaMJLema46mO0iZMOyQ3I
y2bAAoVCIG5wpGqMFQgBU4Siq5mQWOLAeNw5QLHskyGDkFwVsKGF+ev7B2t7DQuY/xUK5SQeYRfu
4RnY7Qi+eEFz/EzGvVKzDqRzP/2sK3A7FKFdb0Dtnp98wJ7A6cjCLZIUHoDwIblSjCf2EaltTJX4
tUGhhpyCWtLjYfs8dqGTJHap+2OX8kqj8tLdOD2FiWjSyIDfGrO5Z9eynZ119WcMWH8QWTV2HErx
sy7hhGP+SKJbnwdMrd9sI3qxhc/O8a6XLjTFOjf5vH1ThZ5qeC/51rNB5/DRWaU0VRwFo/iw0PcD
EIoW8PSqnk5vaO4Y0WeOHzSeB1ORod28nwWyskXn28S5cmi/XYlwcHxX50XD1S8i6A22f3A2WHOS
7KyIpSzV61lvn+TMxXa4xcFxHnnw9miQr1NNrWIj3erjkeZBZgo7J6J8MAQR5WwHiWunAFqj6de9
QTRf9XSnEsDzQrkxVY70WhOY94hhYtTAS+KpNG348DkfNZ6wrWuFHMjHC+hIs43ri/c5Wu0JV8Go
EMYwuqbtjmYSeZh2Y2pDaS+ZvEyVfvgPQDfA1PoduJaaANplLcxhWGOk+L8eq7/mZrHBoQ3XgR+d
6njaVTKyHn+1hsPWegIJ+oaAAd+FCuP60/wTNEdTY8KSXzZyOOgX0TRpw5yxRkmws6OQYx0psGOs
GMsBTRtPQszodBQvhTy9TuvTEmn+KHnsQvteYRQMfYekd/oOTiwyboj4VXHkbTdWAojm0Va65M9P
eGR8Yylwx2XZsGGtKSrEx/DceQvOuWjnuOyRDVw0Tgt+aozxLiA0okq5/ZZql6bm4zDkdNURU+RV
ZoMUBJzcidMPTPL8jsoVNP2QGTnz0zKdmR0AjRHj+Q4s7cfOjsREbgy3ykwvxOQI3UQhI1lPyVzk
NwBd9WGqNelIbeE2/SvdC5MBgHNkJoUxgBNfu4tfAfgFSDO4KGtwLdZaGyWmzY6aKvgBXv9zW6nf
hERhliE4yshoFBWYihev+XRWpO+rIfIuCq1cjfjAG7IpQC2lJ0t6FsbcRpPl4qffoUOct6KVEo2k
Cw1+cwRm9FVZfptgZB1GjUEkrL7+H6myX9iUVA2ENYNVXZ8RoEzC3Cjd0L6fZgPEyywwdQ9Dg/uF
BXg36lFb4ydhiwy4RQdjcezisbKi9msq39ZQm72Nm/s8F5LlHCHN3MokyKeNufC0pc9U8sA5DCZy
q80WMWQ4wY6ZdiDZCE2s3nP8UCJmGBVFLwMJzUs4HgsgwMSvSr5ARKo8rHg172v44oWyfCJ1PdML
wCbAIqlBEWqk0Q05wrNJj0+QbTqgBlWFqHtnSHxV7kIJNsN3GXZXNOqq2MbJ2A2BVTLqnHyt1DUb
EbSRt6Bsr9uFaHvsq5FJth8L1/n9YhUcC2oB84FDQT61xWowZu4i+gq0Q6TuYUlOZBL7ZnWc6Kfp
esPfwRiXTBS83IPogT2fqw1AJbbgSvdkhNI+e65rhlMjsuCcFLrYKq7gbRtrGsKuHiCwOlFMl/mC
oB3J/BaWVgVgj/cIlPx+T/S99A8wMayB0Nc4nLzO+zWrF+nDkQEuAZzRI1qWncTV0B1KryZxDQVx
vlMNCiMz3Mu++DWlVf/So3W1Rjy2AbWTPulJvq1CA2JgxTIdoYzTHySSOM1/uDHWpzhwjS20Owpe
t5tPIjdPaln1gI3CjT83KaiiFXLWDANk/c7gK9gg7smyq8k4HxrrwdxMlv7zj/6g/l2s36UpnmHD
lbaEJY7KL7Rm++Pl3uhwnEgYhA9klKDzPXfSGsdlx+6haX+wWtkgHn62eADyuTU6z9cAgDIU0zqU
RUY0mozv4J3cV4pHphNF4eTLQkBEo4YOkL6WXq7UkT7Z2SyFogBicqP7LqY2se0zn8hTcKDBm0tx
JJeampq8I5TEzexbFW3tRWecHQyTdWOnatCDieds5r/2dBf8JX2ejmvZJrfFlR02jGK4czhsvMPX
ch7FKAO8fDoeAVe3/cHahGbW5AodTb6XHrSQxbVZ/K3Kph2FPl6GHOZ3v7YgMpQGITP0l9xzEfvP
yQ+xiAL9ocI48RDe/sxhjw2ZpgfZZiYtQDpWRc0M5anrBNv+D8eCEXfNbiqOMUPLUogaiwq5DDpZ
kLiSEP8IWZJ+bY+YZYhPZo9uFaMSPpIkLEhO9x6TDeHB3nkz5TpRdZQkj70gK5jFrOCs4GdP9lWM
gM3tIOAlo9bS21lxodMxjXvnct0I044Q7N5Kq9JriQiRTGQ+vRwLqqpenWT7f5jxPBML+UwzOBuy
rXL9mvP6TmxXEHv3ZcIJmHyPEuuIebHUlZO+GBfmwmQWMx30+R5pAuedgc2SZVDAZvlePdIUOWE6
ZLPneTsAlEAvHI+hFMDQ59ivuobbI5frAuCDMaMXDoFXrnAjIlhy0rJuglvuVIS34ZIDXUfkGw2y
8LmQCbvh4sJhlmTtx97hGFq9SMFnQGlETMkDhQuBFxYMz0y5x81BkbxJC/VT2896snVrUxQJAlSr
+TaZmx6in2sRcET/n31nMnR8rAxD9SyiAv6fOHP5jeeqOoRrPi5Oe4lNHimcKh2mQ9EP/hHTqYfx
vVcv7PFmv/vX9j6aFCt6uKEULVo4O8dm1bKqRzgDPEEGaU4/MJll3gfE3P6PCG6RT9S1lEhqxvj4
ejGRTjHFZz4l9q0eLILPv8pwqvkWt7sKwoSczVnmEV5XmBXwZ9Tnmanc6mA/b9q+IX2Ee86vTTMq
yxCpwh/qVc/2YxiM0PA1t0Id6qQBDUPp8F0ynuKMS1IYA09N4d4ccNEvK9vM9YbTOScXS0LGdI7Y
OoWce1jR7/kvfwFQ1cIXv/dKn86SipkkapBPf2aVn5COAecUW+Yup4A+LdaHrz2W3zqb12P1m8P/
PQWr77z2M00oJmEynXzjNJo48NIQEevkvIJ4H/S15GTxLNg4c+Nx++MgxyX8k/hf7TqKFFyv8hME
rTBeX/OiFtKY675Oq26CFXfv4+XaXRosABryAlNeaXDEVY35TUvbkaPE7H02vY5rFC6uPKGi5lQn
PBN4Eo8+Bd7aF7+zRgVaWMGCplkHzLF3/qqwBmvYg9f6oemJdwzuK2nbgz3VSky8XocHMRywrdG2
dSodKUZWaSS93YbsJ5bz8uj20ArXPjxMFXugl4DOfq84OyAfOjCIUq2aR2x9qA08dfth8k22sjdC
rNIZqkBhhsI5j792OhLHSZeeTUhEqsdDKwO4PQl7LulbG8sNRE3mvn7eFUDmJzWad7r96wVWirlW
PvFC5FibbPS5mdK3nFbsK52U268bKntG/Lf7RSxrYtdgi0X+SHwzOgFnU89dJIm3F4smyhQNuKfK
o9BJbAVFHX8zyagi4bh2L2keTp4vscOIBVWtmqgI1bXsX2Kz6tQw1jgtzibagVHMO0tlkehq6lGj
mUdRspwTupPidjXygla3vZRzuS4/PKzWMpqUWAJsf7cIwMUmyFSZ98BerZXYxY//sV4vWpaO6bjG
pppAKhzKxivA4/QNZ3c0wUFCZDdfjwgAqVgtW4Pg1SaKXPbEwB5TNg5gK15RR7shWahGacn7+t5S
f+6V+ErUIWhVZpRpQuTzG0KNgNl2Dqsyzczjs74q9jd12b6e/4p9OOmEWYdY/WyBTAfj2TGPYdq+
LZOFOnrMiwkm3kOS0/4A7VcpbMnGlzDdKt7wzMaKZUWuuYLGY6UeeWzjbh03ol9MfZFZ6WGt6gQK
SISiGSZ/g2rn9V9kocEaHHlK9vO2l0XR1Y/zQDwBHy/C+VnUm5OMU1/nC5CUznAOd6vx3oQpVxF0
tKyG4MpYXFD4dENNIkw+J0+KujEkIH68urH//Pdqq4gb8ZVJlHtqmQHKVUwIK1k6chEwWkwx87Q/
gta48uFHhs4OvNe/ifk+BeFjk4eFOW91Yv0Kq/K314fthdxIbz0HOrPYNB+pcgd7t6lMhsYAfk7U
tuOTrC92X6mckuqQrpaLN2BCUM72Fa3y0eyNPo9/44TqzUXGuWwFU/QQTxYbEjw744dZbK5oqh0M
MlDkVKQi6HNotsle6uVB+6TNOmcjsvD+I9QqKlygqziIQ1bOAWEzigtIzWhL/Mgdj2m5LtVrJV+x
G4K0HknL4tEGY7Y6XQjePASLDBPn1uvqN8QO6AwFhZVTEN4zrupIPC6f6/wxKlV2/TyFU/jzz6qx
PiNXBY+5RtKlfdyxf6ffYS6Kei4wYTL9Uc/FFkYoxCIpyulymjXT8hBA1KoNuIKCkX4eAUUkuIwC
dkrd6bVRpmx70LvZQxp+a6sMaJRqNdB0wnQSr2pTsDFEG6YBfzoz1PGaAJuU9o+siL3jw3bwktKN
MOoj8AS2wkF0eV5Y8TQjoGgep38bIfvW3u7zyeN9vS/QLZsWvkIHp6dmGHWNN1FhqjIWR51ZXMFi
hGWgxa3v7J2rCmDiFKvlv3FTxmt3+JSCYcS1GUvgcA0AOkdNTKAoqmhYri1SF5xb5ti3kL3HLsMx
mFvo9+j2GlMGGTkDsguuEqF/qk+/mWeUlGt316Mjt0NNDYrV7OXS6DXVllcBjf26mBsGvJq0CDHI
1C/soe9MQ8ys6Wsq9TtnmwyMvUxQJCc/LK8aPARL+HUp9yL2UW1V65kCrthn62QfypVqv5rNdzVe
erqJhsITBx8vpTtsE6AJvEjDm8CqbLTIcQPD6s6pV5Xp0/ctjUoOxpGGlyI4a4v02PuAHR1VB3M3
HyFflR6ZX3iDubhTXN0lngufhvgS8FQJ73s5UBaxl0OiQLWBYQdSIHx5Dh863pCVpcDcz015Nttc
W4Xme5Uui+VxX7PmVT/bkD6qYfeptXuep9tiqgymihVkFamby4cRXND4rGeqm8XeKZ63nfVX4Xv2
rS0WLxXQD1eaY0I8S3ttidG5HP9fMlZWEFtRCXzwqDHIESaKCZq3V9f6eTUbGwZbA5tjLHixjop1
Z6/YHEIAwO1tdx0vF2pddm6AKuXdqOBi1cV2xJVK8wcw6ndepM6kM6mGSsKv0D4dVf9XRiYMC8vf
JzwdI9MQaCUnepUSiPP49ELj9hFXeFbInnc4MDn/b8g1X6WXPSvm778jhkn4IKSofJrPB8O0XsZH
vRCY0HIZj5EURJ4A/wtEsXxlJf5n2VROVZY9tkK6v2kP3SOO8LsgHCekG8aA3EPBJb4ir5k4/64n
LGELiiNIYbUAYrX4b5yMQt6D9MQqMJ6lnTLPRGnl7fb327iWZkt/NRF7+eEGb07UOILXAvp5KUKn
EdYzFcYn9+SUGh0zPWoKWMwoKeN/I7Z8ycRezCV+xI4iPyBDAFUwrS7SQL3WEm0LWk78uaRFwk6N
oN+EX2PgJcNBZ7DhtsV92XJRncdomV7fS2YWZ7aRqtACOf/wTffQirVU+6ViTZITa1++qvLJfn4a
skYlnkecxiqSvzeyEN29KiVUF+w0Key+Lzkf7NFeMOHTbbvnmp8ZaRujxdolwnaL1YFyAc38ciHG
Ex+CxYMX+CKPanik7oE1WmKobIFCU0pQ4Ila05j0/YwcgImgPGN8Lv3iGhvK1jyY96dm2Be86L+8
0j4/w5pyM3aXPEUbZMYFMOn4OC+z2pgQSLYLt6cAlIG2BK8K0MW6AgATzKd02doTKNAlKwNimp/I
iy1s3fL8BtUMbUqtQV5lMti5OhbuXNUBzgH8X5Qoz6AY1V48eSS/ZG6/cXng0RoF1cPB9S2oXm4M
SYNyLOoUphy23XMqtRAAJJWNDEIRBZByZlykMNvNR6eFXxuf6wBXx+ASo4tjSj470COrkkKCKVoY
ZQmnQighRUacj8V6mNjPO4caNyxAkpOnws4Xmv9b60cB/4KV3Vb3wHnp6ZcgZCIALG0A8gincJkD
dSCFz44Vyk7gTE1s1Li2bo3vUrca99dZj86A/weUoOhwRpLwjnvjvCWbBscCxgRYV3axp0jV/pXz
RfNjohJ+qcU4a/ybGh6o0sMZgA9HgXeUrF7GHYQcLoPXCJw1u0GwJNrDvACt+6ezkyIPvY5c1VrR
E7IGPJMWQ2G0+alvAk2IBqQkE0bVX60lModr0AiKvb62wvAsCLdOeO/xnBfdyXRxDa7YpUgzbCCi
rAYPb+AgZtETx9IPaJyLB8iZeaP05h9DuJzRjveootr5lyIeDALgDkO665bIgkqw+eJOU5MnpRcV
XtuFk8g1JHOJqXNO2SXxQF+K6sYDjFtNdVbcW2djYJ/qRE5ZOPlRTdRdI2Bb8/3gwsuraDPAxKGs
ckHx6C0IJDYgGvL7UXYDU6ZECP/5fVIvxWQ7BZ8K6L6mqZKGOhJn7tG5m6dWRNMiPZ/8mbBXkzzo
yg+o0/EUy67OnLOubfrDWjyxUUezcPBHCnbZsQpAXlVx+VPUGomJdDw0cuc7Twr21WySTyiDTeN4
/nYlcRjdwEC9F+Ve0JxHoyWcZ4xvR7b/RwN7sJ0PO5raOG8ZkR5z3Qt+rkP60NVYeyDUdljLKkKi
7f9uXDezHE7l47xKdLDMN2cdlO1Wwqnj9iKiYz7SYNtetJqjQgyMFGnVZFsbHh03d9xcQAh3mhZR
YfDPwYcl/BVyb92TlFu0WeD6Nkxr5Z9MFWYCpmDsb4OEG9+vKkXhB3NXpKqXcrrhq0+kIP/1LMtV
Mi0nxLKBqCKubjtSZWi4PobaopwHtVgbN1oTjtwAdQ7Du3O9fTEH7+pgk5xubrMGQgw1YoTJXpZI
TfMJ1cahI0izx7r8t+pxEN1pSBkEXDUjA1IkgkoCgv0A/P6yTTf/3KppGROauGWSsI03gYIDz1DF
a6vJgLtkSs95kG1NOYehLgbBeeUhJXSO3sSegR3zYo01JKJgJ57/8XuFAWv9CDkjjzbfXizCB/80
nHiI2LFi+q9XnhrhpYOVyBXq2gtIUQThzmWBiilg7bVWZlLttC8pXvH9m4evZ879NR8L6uEedaKd
12+6Bce7GTX2AMZWxivme7oJU3/9vvSuzEptKzeQxzZwbLp6Ntjt8X/Vn6Hb0n4Sc5CPTOmZy3Q6
1kks9wEBx2Qn9yEoVIuWuJl4nPuo3gRpCOfzuWHIkqMUyL+Tb44Rn9pteEI3qlPG8wLKsFAIBOwH
yHTTQe5yMlcLSztq+5I272iaziJf6/AeFOL0A5YY69Mx9Kfevao6S7SgRiqv05C4ZWk4wcGmp0Jc
YEq2xRfXN+BlbGXikr4L/OvjLi04uEc+4GeOank4BC9Y0tfZxkLcwje3KArYOGuZ/aaHse2Vs7Wk
swoY/8oLAnHLuJChvFU93C6ocqbu/XiW2MV/JX02BwIC+dcAZ6rY6E+rdSG7yVbLigXfVglDxZV4
p/iru0Lt0Yh8GEdmgxjStbBLqIdfwE6CloFwilyPIr29TEaCpsVGkIHUn1q7UPot1M3dpcTh2CqZ
4num0L8hRgOgp6wKaS88PrSOEMuIpREFzG40OBUWg+8mODBgYPcPTJb9ajbkcfIowh/sB+gFwtAf
UNZHM9tpPmVfF6bHwkosFvjDYnuzZOPg/UvkJNXsyUqzGBOa141W9aN5mH8yNy7oClQ6MiQXHVI6
65sM7JLtNtJiF2rkbKUKyW1ygCcTkh89e9hMETvNtS8Mc5ZV+iO2Fm35dmC2a0MuOo3TI46DXa7K
UEuymghwbWiYSrB6Lp5QTc0ddwdLdSaEkqZkywxFY88ZU/Usu9CP3D/Q3M7YYnemznjZ/U+CgVog
yoB7Hev4XZB3lMzuA7oTUP3H8jvlEdrxyA3R5Ep3+Jur6Hxc5KiBFtUkuJ+gTcQX/cCZhFhzeZZF
vpZImbLNUCK7/NJCGP4XceDmSxhnFZ2vo2XIiwIoJC+2QdYXnuPeSEgqFR/5k11R9T8qIR6dgaqD
awn6AFcz0szP1g297b7DWcSAJZhYvEwgwglivYw8QgOzd54slaFP/+JfFZHgq1Q9gg/QL1N6GwQ5
QeSPbimndRKiMWgYok1nXdBwfmHSdlfeUe0L2RxXrvaqu/atq4amJLkNPI+GqDsFFWZWiARwVVta
hpIBfaAvJUxYl/gOVV6uQgv2UCQPhipNhecV5c+mEVYRgOxIcDrBDrpP+vfS1+rxGddujOjXzD/R
iqRKyuFYVfqu/IavoBrkKyT3OZmyoZGrgpqzxmkf+2SPHvzk87Wteorj/mh/6kHpFxVcgRDIBNxw
jfPoK0S7Lubnt57UQcOAoQc3w1EVi3a/Pehjy8GFzUsIYcYmnlASerqhR4a/w2BEnW/kMnfSHQED
X9cgZWl2y30/72g7SrZ4uCGUwZjjpcA29PM+X0nXXGBKt/0kH3LCm56JqL6p0+9+iWgZw0J2zovr
hx3WAHWonvMl8ytw+QfCf6+TpzOYSEq/hL0BlShEvOiiSOdTB9oExGrWmw3MNoWJJWUk645y5TFO
sfa4ktNHsV/alrp5/K5V4hYb5G2Gq5RZU28J2gdFFzjNdNd9C2J5oxyM8cHc4f7YoJtOpIHF7b1F
s4YZzSAJkdyfGC1CIBORMEDacCMa7GQkIddjk47d60+lSwNtTXy7h31BFoAypA8MUSlsZteXJ/83
a2bDszvb+H8QnVrEL2j5nmwr8y7bez9uCHZXITD4V5LkaDe4Ry+dIik/HAddMMjTqAC9MEoyyxsS
g5At2VpYmMnRbNxN0r7xlGu2i2gR0JX4cBuw4ozuDvSFHA9xLi6STQjBwyMGNOwdHtGFMfMBeX+k
1D5e1/wd0InIxvADHy4zlRom6p2LXfUh0BroLIm+6ApiOj1KiJjaqkfMmQOqMhhI6xRQ8au9J+ed
3Y/9agRNnB+tdfMDBeW8cnWoTxpORF0mRabpdoFnipIYc3XYNi4iGcYbJVYHYbndRKkjfEoYYI7z
WKhmhbqRHmb/SYd6z6nw8kKEkUaISJM/th5fofhNoZg4iuetOxDUREpsG35rqCbHge4ItOe5pU0A
RqKJAbE0xBMWR8nFXvqW49ItT4ik0Qvkl8Ev9z8SEPerEjhrnuBS/iax1tawRNRjIU8JLCjgg8vR
RAslpaPjuEurAxW3hsPjg2bkhetX7ociNLbHjHJ7qagjC3kRVutkpIm2KZrmBoa8kIjla9KYWRMs
UtL32sXJsqRfUww6f5yJTHEzvHTNNSzJvS5U8f++mBT8Xi1TmRcDgf+HPObpHPPa9nUDYVJPf0GH
r7PwEcuUvssjsPzKLT9htGxC9SsrKfM8dEFPsfLSvnFZhsCR6TdUqLCr3mIawXsWCwwwnET5WmfT
MKwYT0T+vM5J6LmmSBHlXd4U4FyWp48wfzuCoOKIir8aCJi7kUJ9ukyW4IN/fqS/E3ElrUDY5q5y
SfRmsQLojrJtZMhMnaPUgIyeTZrIM0kMkxctFQJ4CMVz3X6F5vLtQIrv/Tjw3cKu8a42RRnpZugY
1ZR0ZxnBVSzZQ+lNqJtIGdNaFQ9aJBdrjoYxWVQowubiJjTFPAkfzDDPHKPM4iixYInMBw14Ne4x
KNJjL6DWhQXes0XshkG/0onTzuwbammEMVGRuFVjimINMJ5vtBmRRG9VmEuZXhpJ1DUXM3qLO1ta
JxqE+E5WsCelY6wr7Q1rBzFIJGoaMFgFubNBHpEnC8svwY52uEF0vk8/55LaEtV2+RsQn6t1PHYD
pB6W0q3zcXwbpq1TNYLwkczuk3Z+QxjGclotJfbeY655qqnnihLl3y6IIhVEOUy2ilFcE96IGrK8
WowLNlwZvYr9QLK4GMcanIWeed7jCWP9hn6U+ibEdcE1vprWP4HsRzxmie8HoNI0uKLsPVRJOgs8
QgasnPmYoIBm6ShDuedYsE7e8a2Jr+4gMznFhCnjRmS/h6uIxIlqkGdVij6hCzKVBoZNXaNQZv2s
YoMFxlHrl6EzmNrtS4R0pTIh4nv4B1Awz9rlC2c6mJOmUB/kQ0OlqnJSKKerMtvcAOt8O32cZf9I
pc5QhSc726zMyfWJU2a7sYTGBAN13+z0YdhlHdFDw/a1Mcb6/Brim7ogqJImQjtah7TwHOxrDL7s
yH/2d9R03/tUY/G7ufB/k70z2Hnofty/R3778Ta4Qj+OzuzuaTtZV4PROfTRV5zOcDbs+8hTUq57
oOt/cj5aRLtXLPCS/Oox7k2rWHMWwy8UqGgTEb8KP56cM+7xZkRH+V7WMZlwg4HRAHMdYO6/v9xu
MSkXWWkAaWTYaany15/xS2kVCkNLVB7ZwdLELWqMd+js/23cT84kbQzxXY9sO7W3I8feQtarJo3i
s3AAbZ6QFPbgo1DoBGJM9EHATqWd2Tpb0pfREOb9Q6+CN1GPca2q4GB26mw6kKpzoxDAR8ZahdXN
djN3JfldotcTcpVmBsKpWBH4dY8ov8xyNqyotqj/LgzqTa7bD+FPTb5uQ9G+tFeNJY6gQZvUKTyp
5CVm3HL6DqQpiKIxKFncpsgE1oDQTSvBbptNpBFgnZ2y6PY1Gc3wg1trHNzNrEyVrasFZENJoH6k
lw9t3+7u2XGpXaIhgcxApbbvYpHUdYVLjT4vlQliPNg5e6XSHUDXEa+q+95Fi1s0Wvl1UPARqrz5
S/wXV6rDhERZNgfu5iWGpNq8phRvt2QQ3EVgMU3IHcjFQS6+sNVhGp2oNnnEECnnQQP03mXBpIob
PqOBt+O+ZTOvZWQG4Zlg0FL0aRxIurZutV1tN0t07O43wWuveqB+oWPD64hFvO5IzdfDmluXWbjz
5eiasBl63czFQb47TC9xYqJr4OD2k4r4lM8kR8Bx5gwWh0szNkfnEd0ScBRd6WnMU2xY1fHPcZlP
oiNjRe6B1IbJoCIZf+dVgcX97voU88lRfzdlGvciSCeH14Afb2k+7cfIvLMW9tGGqxtMXq0FFave
HIUjJq6m69SCN787hEn/SfQVzEdFN92zV87+sVig05D8njNEWDjsuwGveyAyasAgYeyqxm1/8wQq
NmAxZRq+E0z7T0vE0GECAVZTikssSCQyk1Noy29wnzRV84AvbS5JCqT/q0CL722jE0VzOkYYzuLN
j2kNVwPv8MX4vsssR7Y6wkWld9X73ZCf1NiBb2cstctnKVChQkI8JNgViel5EgxlzwKEd0MKkUnm
NUJ2p0gRw+goI/HI2Up8A8uGDVYFLQvQbRZJxHM8asjrLY6f6h6720z5WxVUaita+A1WTAOVSgv8
JGenLIkTg8s30EvgAu4EAGRcfULHWs65jwG061EfgDD3ZAI7X9dnL0yJXUFhxJ0ejCnLXUnCaLQx
sN8HZqvWK7ru4b/dSnElSejCcMev1I9zHV6xKhV9Tyr/jRoPgpw9y7u59j67L2/J6484l/D/Wn+o
od/AcGn1v9YyAAJ2q4bWQViR3JP4O5eDvoVI0V42EQouNl4xqOfFeE54bKd6y9rVeyELdZOvZIC7
Zh1v7rx4Xnj3UR9CTeJfO57xYtu9Q3BZMy5uNx5bbbR55idjlAuZferOr6OyVt2fLC4+ug018kV9
ufkz0F/mQgnPfBM/haJJ3SGQAqQNF1/xYP4h3cHv//Yo0u5fc7jIuov+SU0rvMUnSrLxfn70NsI4
9RUc0Hictqi31ZydWPviBGm6QMtwLX0oHSNxNZhy+v+BdHWrMKAKlmltCMAdiVoDJv23zN8EGAC8
SKcwmz9PvbHVJlNK1Jc8+82PH6aN8+2dhwj3ceK9ZPcQZXZEQlTMCun2nX0xM0JfxkBpSoFHwz57
7erY09rFHqCIz93sGYPsM1XZi6p6alDfJJvHVdaMI9TL1rv6fsL+mqKt+OK/SVubFf46i+Hf76mr
pyP4LsIzaBXt1ikvBc5WiiWKJBKLuGC8CjkE5rhZ+RJ+yo+JTFgMyuzNLwJn6NfpDMgxVsDRRCLB
nsw05D8E3nRjltGEA4t9ey21UF+dNHuwpIIJ1tdc3t9mRay7Qu67ofmb2tfJr7tCjDu1ZwB3Cv+x
Q/iqdTrsdwslAGo5hVjS56rPD5YM5TxDeSD2aepXSO9W1SHJeL8/vmCG+aKYtGzZa6Cz+blkYVF4
1ErNy+kXG4LHrgcoLcYv9eeobq2fhDIzlqwLOupX7Ue9rCTO+g0uB7qGjLUblpLNgInh5DuvrR3R
aq/fCeUBUMRC6IgTz+e3BuXOeiz5aQ+X+h1/vaoKVSfUTAZKYKomHsyKp1QETfrX09hpzu3FWkiZ
g6tIsatZiQwfp+v0SdVUHbW2dbwA8NHVGEfEt66SgEujV3ItG9aBsKy5mY7KHx7OK1Mt3oXLnW17
bKKor1FtOE8etAFhN8MiuLVL32SBLGKaJlf4ZyhQOvBJuIatyPqL1w29kR3smldaPqcdGMHo/UP0
6ORmFMdNkIgNOFT0zFmM3NCaGK75g7kPdkFirgrIEhnbkbm+Bubr/fKG7NSCPWm9dwQxn3Bdi1ra
UvFj8/tG/5sQFY8Trb0CQkPpH+Mxodu2ilOHOQw+XmWH2TZB9lb+8ByFPpmOiHBSUVBxmi6szdF7
WKxd99p5ZaZelh5dFEgUINMgxdXrv5OOddEe/rUu0Xb0Mp9cnnskzp6UELldZ04fNRd8b7uvI+Gu
kaV80VRvAQZbTfxSrwv6MvA+kxJ3altosby+dlK2D967TZkWxXsD2I8RV2A4lxCaDOqGQpDpH5xT
L52UZotsswxuJxHFl9+gAnVsyDb/aVpYtvxoQuZmaiXhv0ClRxDhKBOCl7C69q7J7cXU1mV3i5x3
XU2OlmH/YfaoQRwSBSj09AyfjAn0s2RETBKKtrt8PPUR6wJgUSWZPTsQQ5DFIp3Cjeh1pX4fcPal
ihV/Xh4UiREGR4xx8IExQ/JgnST5d41TFS29O2mwjjgGBDUxzMwNikyDjdZKaWowpK2VIHpTHy4g
INcISzJuKN1QmeL8+piZXcKQ11nuDGELupCb8zHUlcPc2b1SwF3hVCWdM3r9GCllIBrNDvPbqilk
KzSVQUFmAiGoOCrcr+XcyISyNMke35rtKmtt1Wf9OneNtRZuiJIBeWQR8jg4i+F2jGG3jB5PIKbM
F6wEHh0j7kfmId5elxiOoU4S4qPjMhd1oimL5HyUwi5yv1I14bdxrovi/PwRHxIR6oXQDRk8iZt+
8Cm0y0XinfS/LiB7VuQK3tInFH0Dp8fkv997zh8pHlIJYUexEYQg4jFhhWyZshGMo7ZwdL9mhbva
bOdzDq3ge5jsOb6C7crj/AfBLvHsOFH2CJmJsSpM5hjLio7VwiFS61pvrgyWuJQGH12zpccLDOcn
6YtCtDkd4oG1lHhSzpMX0g5OeowDZ/RaRne2YO9Z723eJ/KZ9ITI6YLb30McOG1Syj5c+9LFMY9B
hmxNYI+iXZZmmIyzNwcyIMdVtBjD+XqY8XDnf1dojkkDD1m2w4j0NUGUFcx09fodRrlLGL7YBSDE
iN1ZeCaH1rvFYZJG1a3rIem3n3G5IK9cSS/qz5h6DdkXd4jMyEo9GzjWxKQcGWCB5W52LrjAEpeX
7GHIh4mEeOKQpjoqIHA3Na308MSDa58W9qWGnHZnzo4YiUJ1MfmvWIGxITtXlFulMoMt2Qgdr+qZ
8QfQACeKmwB/ffeSDvZQrTKwFNaDEJieq/yZVW4+Qi4bYEdK7TbZKMwtyF2JPt6/jcOM5F9DqmwY
az+jmAQ9WiJoJFw1a2x4nc96XuhvpRugRNl2KoT4DVN/9kFyur/COYT4gwjCqkEpftaa31W58+XW
QOvaWGRo/i0M/HEBgXC5SfjIQCBADlQy2MZa6cBeYkDNeTESjJbSWLGtzq7hJwNghFAK48nGTp4e
iu1HzvEFy0xltdPdF0IVm23RbyvHq8kj2Fc0d/EJfHaqFgjaF3PeEzFVfk8fNA9M5RcoFGhBrNFv
2gUKpfVuUTIWTHGAbrMLwgLUL2gnbgKfDkBrJp6ri4I9PRx0lCZzv2wpAH+BAEXT2MrMrpKctrtC
9ELrjobiEoNs3zC5YceQduwrg7aTHrVA4hjgvToVszVwxE+8vmNKMD48ij9r2sHmJNYSkARz346/
28oT+5J5jlq2YfhpbLRyzA/0KpWyTuLdp4hEivD8z4BewcYSkBZFGhbToxb7qADm+gNv+wbdO816
aiaKS+Yr6wHFknwC3TcW3CFWDRH/NrC/TPZSnc6INzJ3CaCBvT/5pMZyUDvxJUKwI702DSVyYrF4
i69VQxav5aZrevon3If97TJIrVhizJL+AaDAwKf0chmn16AgCfF7YO/u6BvisfCMkn/hRUYnrmUK
C2f+64CzaNZ6PLQf6+p0IzxhK1QV6lwncduVTuUxDaPCnNr4ypFbErYhG4fhl0I3DyZsQJaQI7VX
2zPxijRO3urU7dDOPkfsZ0wV/c6AU6DJfTGq9RkRaWSS99TRCD3+t2YhaJuLtrj53pEOUB56rJa+
ycqnMuLVfn6635HrsmdxtTtljZ0MWUKQnkhvx8JxAhF4sh2LcSfS3PiqhjPuwgx1qkIIBuXMAswv
RFFy+7HEfO0TUCkOpx9HtB7usPR864mxKxBpxq8ooH2yTRZstmZulf0A1O6+uKsxhVquGoyG8nGk
ubSi+xBzSAc37Z69RbGEIQSoRnPDnwIxeEgPOlwEGpQ/d8NlcgwK/b0r4jz0HyRaGu5QRYwdI/jK
35KZNTi1Y+eovb9gve6JSSsZG3NrnUXPTnmFagsip4bQZkggdyA0+uDWlUiQnmUf1fUJmBQ3iSNu
IPQM8E3ZrnX/rxI6+EdtGY7g8AzGlaylhG6KDaOuxlRHPaCFUv5JfYOn6VxQrvf6A/ssTo5V17r8
StwjN1VOkFd/ngW/LSya6OV1QfxG8aF59tlSXNwa3kgvAPI4hKxW0q2qdLT21Ma2yEu+cPsrWr4j
TIRVQMUd+WtWFGrAy2CISp9phnaqM+CMrN8XHxyYsnZjYKr8f5qzIhtx23z/dkqiKMB0ZNpq5bfL
cujhTrZv2UM6SFU0GKi1BnPlcSpRFNJDMuBNVnXZnZVNiRBO7Drp7tVLbsgbP+g/fi9MKqAFI5zy
T5HhQaJuAAAr7OZo40YGVeMP+rWryPfh3830DsZfuaKIsBnjTNlg2GTKNlFXhNRgW+TLxiGNhdtd
HJQmWX1gsUU78RHDMMHcvBV581ZjsIkRKCWPV5YTywwMLRRWKgXkranEI+/n8I8vpS7+zqGL1Jj2
Mfk/JPKmCb3vh3PKSaO1Q/WjVwHwI6FXPAwqGlgM611gUc+l8DImxrRlfgA7waDgIXzDExYIKvTB
CnrZKazaWQ7hRsR72GgwzIrvwgTarsoZcDAkBygiWe6GCdUB1Qpy8bZrHKQhFmWVlZUjI1S5Q6MR
c38Bv8cV4tLdfnG8iPy76upHbeET/PI+6yToZnCRL2YLF7DW2s0l+jKN7W0EVsF3tKKQINKKT0SS
MiQE1ZcwBj4OOp/9BtGbe4VbqcCAFFgDqKCOZPCO8EvZ2QHMYJNsPHx0kmM9Sidf81tRdYk1+xvV
jKx9+XMSebK61O+aiCmHZG0MHZ9EmPPoayoqq/rjrO+antvY41DUpqpKzVFHryHJurV+IE4GH6K+
lqz242fVZQ/dYaTFRd1g+9hvP51WvlSBdA2NCrUG8/26/f+DyNOVV8ocEvslbpD2crem8AvaMfn9
Bz223TLXNbWxZ5bF4qDILyCu28pfrmMa5puJu5lXh4ug3HJwbAlvG69q360tiSQas7wk9ZGjwg9m
f0xxrR2ws378IoswLQswolhLipfyE74VvlEXqAjg6RCrDqXaIyn5+e+YJXVownT7PtzrtJ+1GX6c
NwNl8PiEklIEEFRUtfQo44XPMzzMcFlizHhaDZkIBQOj5voYY8txCh82pIZkAT0+90EdMFsfA5qK
bXASoY3bTYloTF6sDh2jiUdo6y0Amp5aOyQePmRpb1ucZTdzW3rg1aGtiIcix0z2TI7jd1b0R6yL
rfNDR65D8wMdkATVmcKAEOweRMU/BD0sLoFGnvTMX/oGF1s14GCSc8VrauZOy4Qn4ur8ETUZ8D0m
qF0W9uFnGjL8M8QZW/iTCma+a4bebCnxjfDtyDH95HOENO2emUTvAOvyfVa2aOeDNAZG/PiPATjV
z/OAB6lTH0RjBhiDoMxI5tpk7x/mXaQOtFeG6Xy1jn7IExiMDeh1rQ2tMQzEU9c/JBpOBOkzDtLo
IJWEkYwjDgVRyjU9qlToGiIFw8De6p3Wq9UIiah9uJ6K9wlXM6zkQC53QUa7FMbKbR80DGFmF+Y3
WTWPc00LifaIUVEZ4IoABC5gdJE0a07CGDHANIwy4uUM6j/yNHO3jGCVWhFPNso3quvi2rdSBy0I
/vKMbaBJLNVhLx3j548Q7Tx9xnQ5sGVXwSBY+LXpOilWDMiRO68yaa9+ov6WAIFeezxOx/91RfP8
NG30sF/+qO5741YMk6rvKyUU7Nb/IpTAPsLwfWcjD0CriABdAa7YHKY7stjPREXQIArFqFpO9lj6
cPSc/7uBaFqxzKLhX6WCHlhL7ZbssojUieBFW8Lft/x3c4V9jD24gPy3W27ofIrQZPrfiLUfNxM4
G1h4sPjBOZvG4PJ03bUUmMr3tEsCzanM4DMrez4RSLXDt+J/pKpOFh9sqv/fUQO+qIEOhrkqitZe
OFdlrtMNd0xnraV+r2UP2s2FrVFvMs4eHRTBBYDLCOnB5ziRwMPykMa2NTsEJ4BI70Wcepo1kWFy
AQX5Sm03zn185jEuJfY4lucdkAvUsEqs0xzeBenEXRnZrlVe/g2rtei705sycjtAf+9hl7/C0FFl
q5Eefvxje4F5yYWX+CX0su9xLlb0ReEMLcInAl24yFu4Ow9QWlKtW8HeNCw4Wy+PSXW7ITiOEZm0
rJS6dy+RuhHScG17PJ3lAGhYMB/F4KYKgWbTv4mN2bwq7BOoYqeP0mGZn7j9iqvFibIzJ9gzti7f
VNFUNJMMFh6PIZdVot7zvzLRfABYgePgIbYm9KeGcWN92Y3Gm31Ohoo9AUGMrRaZUxhtVnsQsPJf
ATkOjN+IcLKdaV/AGAmpxewVonbxFrJNWsEfugo1uLb2YuvV8iqFU79CtHdxlOnmtu0tWUmVVNIF
ZLEb3qgiW6oB+w3rjkLeeFniq7aMGgXRIXwX+JuHvVIVZNqwuyjGh5scZqYqKa0QatWrOq0iuZSx
bnDYbXMV3b7Q0EVSLJ5Pl9mc+2ZNKlplYu5NXwOhP4Q7D/A5PifCCowLc/EBDB4fIDKkIbZa4DEn
v+xvK1uh2N8TVeGaLJ8jfOUwYFKTUiD2w7jDgO2vFgIwKt5HihFVc5lIKVIiY5QeLuViUT3z/sRT
2Gkp70uzLbOueTjTK16GhyHjAja8dnV0C2hFiZBljnT3BiFlLKbegmI38+VWbQrKR58cfKNY/iS8
gNQX9oeSZlGHJFQsWhzA4pJnG+3xnUgX/3yEABrsy5ZjcAEbgyEpeGSKFB8W5YfWlFBO8qvxv8CX
LDRQkfrXan3OflSE8fBBfVf/8B8wSGb/3Ut62vbzbspZGqFqQP6MKZu7Ew9hadO3zX/DbZHdnqaS
MsC0XxA4VFYkze0PE3Ewvxn/5RsgkXietTcXeGf5GSVJt+6hFM2JmIud0QG52JI04kK/9Dptr9ty
2j0VHxYCXtF/YDQaX2bSClY2TBzcSLxLTCe9rqSZPgRUl1gm83aB3BjYxHLzhPnIr/oW3nXRT/CK
MtEifUzl6b+KhuKyrcPtbx/04Pign5mxBfQvGvM0JXmhKceb7IHh3Ab7GJRX1SZpUFISlkXGD2HB
cgb9ST/U3pv5BBlHLOCTWQQnmmyl5KzhRfTm79BOCzbvAlauGU34rzb/Bfx1pGkFkLWmVxW++GFO
DSQjWyvqN+hCoEmDdzCbrvA5+kcQpao0A6/Hnb2DoJKOMqSSNueq9M2OcpR2tg4e4Bg1Z64wUJ5M
91yBYzk1lb544nl81qq/awrsNeJEpUEQoTyJeO63UhO1yrxmHB78MwrDBWBxTJPv5gmWUYY40QJh
ccqwkjMHhEL5Wz+V7AxQSVRpeE8cyRKMxNSTWRIVir/2+W5f8mJ8I117tsmkgoeMwi3T5xVGGyjE
8wQPwEo1Obrqn2/bofwoP1pHb4tfhOdknDCPG5LYhp1f/zMFx5GSex/EoYQr+r7p+EOVmcyLCzDR
VMarcfWWp61msthJ9ncQ8KrJajL5lJJRLRwR2M8g/79yeFQ0asV3lo37CHh67Xm4IrYGc8gWZSRP
RrQJ45V/TbfLnQs7esCMd5OSMbcdIQlCW2hbDG4R8VZPrwnp5q3NOCTaGTzqhDHW7sBvh5TqlCX2
T3fxx6zngJQlELKgGDv01IHBBhg9RPMHeWwK2QkFAQD9JOpyfGjLUX/Pvp6daeR++K0KXD5Pv+yc
H+uZN5YGTEq6EF7PEMqlsaQpMs3bI0RzOf9vScDd2yAbrdILYsKsvk0/GTrvEuET4XC7zuD475DI
caP2DelBbYfkQMVhMRQ00yNROGxGWT3TrdPv94j+zJgbREEpue1ZcYuUk9YMZntKe69YVwvwOCoZ
Glah3W/K4lfFAs4bv5fjWZSopiBcYEjGObBhHep10bmBn3FIXTze85ygFQsDpc13tNdWMugPWQoK
0cinCf03RE0/K5se8Idcw5t8koO3CIYncjv+fL59SFkRbJrrLdrc1RZjneuRl1KWxaNTAPHOkZ/V
VrboR4Oseq2I3HP1/LzmA5zbYCYgrJXO44lEdxMT11IfssaSJnAlstZ2QV5bakG8pZL7I3qf3xvW
SciN10c4u6Z7/t7I2oG7jRCY9oXp3u05YLOf078H6f896/+H91cs4olzjVo1UUQQUlxsJV8sPi52
3lFXx6vGyFhbemtw8C32hFLUe2WI3juNjprc8zfVPbUwFF680OZz6Hf9/bOfXbc/zbPQaZzTCuFH
1akEp6dETA4oWo4JXSi90n0gA74V/GPMnjNBBtopvYD86LkXYCQqdt1/4p09yZugT7GI34il7MNV
zXuxPyD2TpeF2IV841npqeHP0/5oa7yiCErAXenD/ZpyWefthNaDWK1pitI+dgCNDNc9Hfeb0AJI
cvgnLE7+ZQIZgdB9bG9oupSBL1yyZEiXuFMeC/Ul6Z56oVlWEhwt8tXXH1v7umG2COytufT215Eo
7k4/N7W965r/DmtlSdrEfcv/nQ3JTNdp4qjtlylAGCrNa/NT0jaydtZePqV2DnNQAXG2FS7dJPi7
h6/DAEdkCDkoL1cgN8JZmafEFFTF/+UgYU0o1aTQMqOOyVb15TooIt7cr7JL8wzVB+XcmpGPQ9dG
JeGMOemcSKZyN3jXEGrjlkFLc08rCjruDAoaVb41gjAfcz/EptwZ6b1yx9A3mJ4Gnzkb4ud+Pwwm
HAb1cCl9sbdNYDNjxUsWh8B8Ao9QVHFwQ4n7C+mFsiXqwNHRII8ALx/CuIL5kZFXle/jGyym9gSj
Q/6ISt/qwqXZHd30yCh3EV0EgH+tBDLrOKz7Wap+PwuEBE9VPXUj1upmvcM4bmLKOQfqfKW3exp5
rfE+Jgmj0blBwysk+SIAaIREnD5QRe+5B2DeNjq4pHQrT1H3NXBs8BJtm0oQipN+szVJPdkhpdty
YcZ06aCzGaTVmh0ksZ4GPPWOMV/EYds3tEsF6uOnq7otWalUQxtpqlTFbl/x18wm+pZkAYBRdcUh
4UHLuFL3rI7CNvLBx+I6fKcrLsj7O3E+ygmzrwemHlLIk8gbxVL8EPkJdBl0vEkCxxvuNIuu37tf
6HF5Xy9HippbpR4TeMX2tnyu0Fh9Ejqo0YMHs0PGdqo7ZMQqaHEipVMwz4bX3/ggTpBn3hyInIDH
crUyYa0ipthTbIdz/NXMO2dyXPNYp08Ma0y97NJ9+c7NQ82cLBgXQlNESDp7BI3zLTR/xIrdfokp
xj2aW/2TV4sjmM9cK3L1gIqx2xfTcgxw06QzUjOQXiG7OU0p5zIgFnG5ljTlPSDYIzhlIiLzbx8N
bT52d1uGaGZiTI7NgM8ffLFdRYk+vvSzjKkxVelm+6c/UFQyf+UYyzMYOcM4ptrM8bzuxVEtx2/p
3qIsk9R6B3pJox4BLUMFspU2Gy2x/oLGa6aw/s+ngTd2CRWARVF3ZjVVvmrLrqFlxcwp/0Xb4eT5
jPGqrJd0D4H5wwxLdNojaQy8/Jim+L2Rjz+6P/3YC2azfGu5q77TkH/jKovqocyApZoKTX4MFSuq
H/FkMoOwz6N+j4tGomJRstcAd1V0sddJaO6osAHBe+QrOckoHNux1WOv0txp8nCCiofQGAyIN9hM
ECD6gD24ma/5KHGsdPyvsJcoIFutSmQzmCpywYuqsiN78EQqQo9z7OrR/BmjxwYvsjqcatRGt2uV
X+2DERLWI9RmvSuNfDunlTetY5H1l4RnvKkd3lgs+05ev1tDVURUi+HhkulodRCoj67YhSkaSb+8
Bz9A8GC34BxouxiWGXCdvW5ZBKmZj4uVZGD6Ltoang6+xzl7ufTlkFKVCzYddCkKPxIQHCG7MY/1
PqmsIjY79RwoKnevpPNrreJzujvvqr+JeuYSuQoEHB0KNGoqe8Sokzk4LzSfXCG3pPOdxoTdQ58y
KeKgYNCizUB+bATUcBjDkIqc6uIYsi//wARkvBwLeLMzY6rx6oiN2Hd7OdKa4X8Mt5ibTZixFVNx
EWgTVd70cPc9BhbLvuYcabgVOylQw4nncyDOZpfGTUbHOZBPIb1uG+X1Vr/Qtr5KSDxwe6J8vkKp
QhFIlMI0uCjLbFVTkpsfqREfvNlYpCMqrFx3QAMIGXh//PewlHFQN52E6/KmVkIrATP8LtWD/uxn
xvSZSfZuIMwHOClQyL4SOUECKC9ReMLuobsEl0r+Nj6vMPTRhY5v0UWGn/kANY/HVoTs5hI4m3x6
xnY5MzrmVsMjkuZOw1SpcrJqu7PUgQevc81eTr3ewSw452ZHqvoNVijWugGTQT0lNFWNaSdKgHfU
f5WEn39yj7wIPSQYSHxAiwyqXxi0D6R9wvtTO/ujatP6c1Ags1l8Qa8oOD/fDF1DZkoXWgQejeHj
sNr+gre8rxzmZLvMuAGrig7gFn0YPs6his2IFH+KHGx3cP77wHxNc3KqL7KuD3wRhTsgBxo07XEz
EiJwh9p+yGHFZiXhR5C/BVTDs5e5uFWHL5RA/MMLV+N4JdG9/LBB0JkJudaQay8Gugf1hupZMYdw
h61UZb0nveqYQBQLfTygx6TKMGx12QdpCIrJFIm6bJldes8t2dYkGkyWV5PQ0G7oLcFTPXOeCnhQ
gMr/LFbAzh2quj8aufBNEWhqTjPG18tK1/9tzv5HiZzLso9D26imHWlObjL1Lncx1Fr6EPeeCloH
eE0Am14kHBEp3goSm4PP8jAdzF9i1FhoEkwgLZw7N0Bb9hDRsC0/p6i4fZ6Z7rLDQOnpeNlM4V4w
fy+0kjKf+QY2+UMRSj4Uu72vSxqHSLc4ebmIxTlIWFkRIlzVpo8sPmGUAcvgJYjSYRd4LxXTNW1S
CS2cNkJNjgdhucU/UxeAYghS/r6M9pOXrLrgNXPzgIEOAAJcmxt2Lr5T19FfkpY4XKMy2GviZwrn
jOpR346gPc4go6SCwygyZ4dotxqMnEoVJtsB5UEL30IdjnbIo0slSWASz+VFvqSxWjQ+/zGQX0mX
93eQIAKJvkuV8Gk8/GkPP9SbND6URSHOJIx5CC4Q1YZz/sMgt5P1n94zM1T8nj1YuN69bBpSREki
5tETet0AYtwrONgglfdPBWoDnvzRWYan0CfNAzCC3QzkhOhWQcnd23OKptQu/eEa1G8CBcYiH29a
LTiyK02tD3+l0I/XLf43+heWHoWdCcoXX6zgbW6LTkt7/6h++7ztuiu8RHT2vZtz8UljHae3IYuQ
zMEjLSDZ3sb0F+X964Pvp7SYX/WabcJTOBWTEUOSlEpVVyRbysipl28sov2my3bnUNnSLAiWc8aW
djysKbQUCFRkuoPEn3FUsdlbsJZXgrjuLhPdFKZ0vcO0P1LBoft3LUgcILLeFzFIIy3HImG00CqO
OHwdd7f1tW1vqCx3LIgnxRnqQxUH0ywtzEimyr7pfvmiTKnq6csP0Pd1jvP36tCXSPjy7SyY09Pp
FYY+83CKcFzX8klDcInLO0piupyqTHo6NFrbjvbnjPuc8/aYN+5rbU/btpXZamxETKmkhFhfWEei
km9Q/m46W+N/BQQvPev9NXkICPd5XYc4zm9l6tRglBQ+eLFWo6K3KFkiQFaJoG29hViaQBx1ehcX
LLuk1gZtLu1cOzs9SSZKCxFiAOrSPluxUz5KrD6NY8pDurgP/yCTi7A2xED4uNqEK+oh97mp4fO+
ZJtD8j6RUh1XVQ/AqTyAXfi7fgQaPa9UkWsYo+tiOcLf290f1WFnsEuGTDBrTiMn58myahqiB2GP
CjO/6asZtiO/i/CRf6XW5+SdZm/8TwIYzx1r1KDnQtmB91/zU1C78gyEr/iOuuAnRraeD+R575/3
g8/C2hLLFk5qDZE1KO5imSxyZw6StSH2Xfadax1sj/Ofj1S9N0Cdz1ivWyujDrpnbF00hTCb9+T/
nAk2CItqu7GC5Opu6neSFJHwbkDNqOtqjXAUP9OggTtgBydBnCgHYgmtonQNUUZtfxVZxOVCuaOx
CZbeXpJz9QoNSKZ0qg49MynXTz1SyPIT7znP2MEVCfcyF0buC3A2ds8mcB/YvJvc6dLxoxlIM+7u
9ELpsEL9iVaFqc69N44aWsC209+HqzSt1a0jU8bqoSZYatsS46bG5HSKuEencT5MjreB4HCGudTQ
l41mLllGBlZ1uCbDCJnlLDUSAUSYizbLETBYPfaopOtZ85S7dfKjnW1GhzGLg0GwGXfxnKPCrLw8
hrxX7MyVSPU4KinoCoRX2qlwJWSv9fsQ+Om7tamQbuFhd9OOZlAlOWiKvr51Rt0jZBmTGDi/xorc
5uIrO8xO5IYknvUtG5rAUdnHVP+8o+mxKWepW5vaJpjVbb5y0G2avMSjZxph8PrLZumGAkXwAsbN
D0qTrXgFwuAnosJDgQPcN7eJ3eokpr1pzPSlGmuojD2+t969zzsmpgAXYFJ4wJcDrKA+5fjhqaFM
8KLGmlntofz50RghB8NkD6DpnX5+x3gMbVlbrj4Kas2gRu1qpPbXONA1TXngRe8MAyvrQCftfKDW
1DWmdbhbgGfpcfePvHtKpoZTBf7eGFHr/QOo5T+7W+sN6BrKrevj0T9i7dUVMFyBKk+zmOZD7MNe
JI/dujoHb93noRF4XT+CbgMZj/dhixDLdv9D/HNps3ceg1pL5yF/myGTjzAEiQ12ZM/8jhoMuvED
khOAXYYPDS3yEYsORjuwkQptOYr5PhmL3Kh5pv7q3uW3CHjzami7MP3/qGGXVeJ7uX/AnW9BgHXw
coEh26j548YdEQ80F2UF9Hff5BfFE5P6y1s9bAs/scFMHv8mfWYwjFGZe+rVMtjwO8Y72V7qR+Op
ygvLnXZCB+F8XTWfgA9Ac2GaEDARWla72u6dldHPF1xxymC5IEGPoaxxyDgmlPmOP98pARCXqksG
SBmyibOwdZJ7na/Dy50egSZn5N8A5BN3whpO/suDQdN+eYPPRX9gxjbHhCR+H80YE0BemfH1C5k1
CQ4llZ2O3mkK1ioRSlWyWJinPhm0X4xP3Iz3yFWZIRkOzYnYGlhufQj5CJyfQnG9c3z8fsx/+QpS
JSoxmjZcXGKrO8lB+Uz/39AFcDdLaXp4WPqaAJy8/ESMD5sBIJhEa/xg5civnQOTJdzyTzUrZnHG
5bOoHujSEGWX39qxKnzkNSiKONb1coP2QWd44sqoQ/yJ4gLILZPdiTDfKFohZ4vIl87WVEswSZQz
HXj3WWNCiJykd0qDiSeaXSBUWgibi29Ma6IjNwIJUT9Azm+4yefNeL4YbdZ4c6xNH1uLlVq8zNwa
OpIHQ5WzEZlWngSgFMbCkUZL3fq2G/iHlAbxFvDq7JublOuT4iCRYD8Hk7vMjDTFIOFrKijsJ1mN
ONgW2PiE34AxyUQW6FR6nz7eyldnrv1vv/hhMJW0veGKn6dCd+Dzy+f8BQ3V6DZCq6mV2KpRftfX
QDAUxI+aq8REYQMS5Jib0NSrhIqFPEouZyq89uPZn2gVq7vOhMcn70dkmAgUbuvn8SeoZV9WQdCP
NLahgarJ/xtLBD4Umi8ORwGh6gIvC7V7ZdBpMkRYx83f4a+Q9s1MalftJwSha/oWX/j7NiBTjN3K
oLa9atCJ+6a4KfleI+Xk1ZJT2N5kyK90Go0hvgKsmXt8oyoFb5k9OhHuF0JmE0vEfCsWFcpIX+ty
FZCbGT5RvZK9UzQpSuvS5mECdtxVOEw5Za4Ti1rcaX6Mr5M8Mttvezu/qLn+dtJCvt9lC9S8KR63
/PWKA+grSQIzC8Zg/nv2eoCaJj56YRJdgUI9ny2Nr6APmdz1S7/aIrtkeU8IpBObrSCxRq+h8pgI
2Ea19KUTsP3NZ1BIKh6E8jr6ga5YXM08yX6hIZyIaC1bXhW+PIDKZc+/hlBSfdBIsBq0VHZZCwWd
TkuLx7DTekXq4X/jjfNVRunwyNNKOfYNfb49ADRh87BieDKKaYMWKx1MhbhH5e3d8Ug3ENtBx5Ui
mJmyGDxtSNZpJ4CF6oARJ0Gkms6kiGkcYjLvYgyngY88J7xoCeohDMO9FL628Zgon0OAyrF37GSi
aXdpePLRmFEJaOujNugOE0z6LQJk0cocubRnmk/KIGq2xfsSSYkebMyZVvqckPmdf8lcmRy19yr1
Y5BAKl6blI4jix5EqSljihsRWFluv6SoqkUxzOtyqRX6VeALejC2q/kXwWDd/zYK4g0NFvXJjksl
QZoAkICkC70L1JXb6zXBFNxVjkK4XHrzWhXq4fwAIFHbDG4Ke1O9GgC1k9Lyy2puVb6jGALhsO1l
1RpxEsJe2WE0P2ZHEr/PwcvUhg43XS93hQsx+Y/594aEYAwIBkCf7ShUG/aLWHOtEiAhSeqRnFsN
NQ9as8/ZWS758hZN5Y8pImTGNZvmuaI7AIUJ+bDkZ9OdNLaDBlwau0y2qcumnv6fWt+h/CfmDXAp
jQVKZabAqWrMLF9OnS6JuYfOYrlyFr1wY/XFh6j6iNUES0KNMgm1MigOt9B5DIfdbTtntuL1UrE3
R106RQCJm9UxUJPwsiypgkXL71JQhGFYud4LPJqMczKE7mL/7sQ4nHmBRRpXMS8/JNJC6V57mhup
KhLP6FBJICRsGxczg6a1jwrn83/vbbGIVhIy/WbSzyexmjbGuPEHzHpvConZxIFGZxyEkj3snLMz
fD0qiGchyJ18J/arB/xcQmlNbKu/BZoI2BZ36BWBjbjLYOsT3e1BkWC+D0NsPk60ursnUJ3Lmpt+
yff3hjipQQrMsTEQJycnl/ztT+qEelkXGmdgbAk12QiJVPVqBbjORJTS9TUFsK6x0lyNHtOW7l/n
FstaOG2w/apMknJuAgJWG8e1dP6j/Iab1BNJVBilHWgZ/MPErX290a1solIOERg5WzMH59a0C7Dp
U/BvJjIok9mNliD+dgzmTrRwRFI/P8KnRXTUcGw/88S1SAxDyP2gIDk7lVInLmjJSQDwctZcKfVV
c2XadqePu/97zcxG1l9/Ub/FFSmtoKdWzK/qPy34MEWB1whf/JgvOo3Qcw+1ZKNws0vyCI3DAwD5
gDg2/SW5dNmJjS9UgiKodU8WZRMWsJ7Fz9ZU368QR7DzXkw0KsTpDYooKxvC4ZAI7ZYhHCkzPnaQ
gE86nHFTKgk4BH0xAQl6PCB2UFway5LzxrcF5pCmB2Ddyz1JYsccJ9a8QQPEjNGJShGpx+sD0f6c
EEJITISAZYLyYaMV+Izo6sagxX0Nqa+iEIC5szUaeTuLc+lYkiQjBI2KS4RfCiNpCZuwUZgiMApw
jW4+fJiIK42ORvEv4BAnILuUs+JgD5ds7cy8L0O5s7/wgi4Br0vEBfBk9Sn53VQUsb4q8DvQkM+i
szS7qM51oTPY1slU0H96S0eiWI+nxpxi36LKp3bKhcTFrVaFeteH6nbDQ+j6SNvi8xEppwVcZVrH
cdy9A/hfnBkWqJbHU7zx7HdH6XvJVRsfYua7xnt5DIkYCvI6afXYee3LpcdCc1AMHpufZYiArUc1
b/0dFoaPuB8Nox0hMKJ8z+qx3OUvvlYlxgcnKbl6y1t8ZrZBKY43DT6LEbK+I4/zcZVh3Y38CAqK
ugziD3rPioIjrFyoZ60zlMfhaf+Momqt0KL0D31vpbpArNXbiyyzQNpeH8Jq1wtQOIhhR6i2JkoV
YCgopJK8rNoW6uFSwxDS39s2/CiixdQK+I2CHbi/5bSwFiyaSVSt0l5MMB1jpFNacQ0JpEcIlGfa
lLgovt8wtZevw9EifuwAKEgXConFqoxrtrX3r478VwnPlaE+Ec0mKMu4qxjNcJeh7aiW1zXojMHw
D5rYaFRuP0BoMMNvxn/KADLfGB9hnFnOQqGa2N+mIsNXli1FblHTYGCF7ffa37lO5ObM5n8ohdzL
6gNeQR1zLvaYDZ66uP3NQw5G48O9e6sT2vDYzIG07z8TaysZMlGsyjKZKq22DvgW7GDA/v4zfvoh
e3HZNq9Mhgw6iuWNm/FuCUXSWGjtNho5vJ5E6ZDxBIKs/kFkeB2AmZierdjxvFpcnzisBVhGGgdd
zQwkX7AQmB38Oh3298FJlFgcMUb03R74iTF5K+5np3EsBOcpJd4AK1O6bqF6CzvCH9/Ke8ERyEvB
niUU+OyTSLufBRyeUbZakuCE8DMMLc+ZLDUuluneE81NCeoICC8sAYjiyq4MkXnbmcvO1DDCV8f0
vzt+TUDAfe73EvvbyMd1wqjwc2kgs/hKFWVmLSSHfFs5O4W/vezd6nPwkB/Op1Y6Wd71xmeoTOu4
QWKf3K7Np/ez03Q1MhYyoy/BtOBT5kFtsSCQ1TKyX1Cb19ZRYEZB8QsoasDSAEl3EGExnEEXyv7Y
SrDij6bcXuCBCjGwHZiEOD8qXVL0HChxEIW0o/DO+OK4N+6lKp9TzoLi2uV8QKaVeGJ95AFLKmFr
Fg0zRvuZjR2WnfhgksjIYiRoW1ouMABL7UnPK+E856CRndIMa6oBVOwblUwk83lV3PG3O2fiL9q7
yXL6ISwQdgZHDI4IKtOFb/pa9xNJoIoqBKq4WSAs0nqOPRjOLPEIILSBcSZTOLSs9iFxLAWM72wY
o8FilLIpfBMe5+9Ewdsf7bMvMqDURUk1AHU/RuxgLiaRos8knckbdgzzaV7M5aPBEznGNu3G2yOs
/HtLiSjtp0300I5IMsTSid7tn2QuHdDAQ+VGmz5VKExkaOFqOZ4z6idXtNsu47pdSJNUp9a7fODr
FOrtXYvTzDNZ8mR+RAmpwpwGHdSjbNg5F6FkpOeswbTI/PmL1kH/b9l6L7xhXtXhJAR7GZP89PFt
oN910pFffRh7owrd+5WA3/hPjULObE7La27V/XN/vNpITIq8VIxyJFNWmksfdMq198cZsHoZo20o
X8cHx/WfoQhs2nqgpqZM2rB9pzg58bzt9aGM1kWAJUugYV6pu0bmHMnzlhA9WYxL9DGknNF5oXk4
mlxlD1U4GrlNMN10AMo7zpgfE3AgbVRAbKHk3mhFfKb4XsiwmuaDhBLqIVA/avqWOAbTT7szRZ63
G8RLJQgSYmpK9YxaZayw9B8GmXUrY7YglF4gTeYQlX67X1GFVyYnSXRGC8SfopUsRpRf4siSZsa/
1MyxoqZuvwgZ4nyvLGZ0F/8qqGGirA6k2gfWUK6hXQ8kapdG1WT0aAonBnRjN7Q7537j/rPezZmA
V24cx1HmAybwXUvloi8LYziZO9QlQO0lp2LHJBXrDuOR8A/GfAB4L0XO1NB5ytqYPhOa7Pyo38u4
R63Kirr9S3asKz9z4zADM0wqDdyXbeB/Yms2+OF3yG7Ao6sa7Dr63ZcHIzAhGR0unJLwvkwvXNrw
dfvp8oemjgCe43RXFKmzHEKrzPYMVMGD28gkPdNXSX8fLJM8gwoK6z59cZi0RUiyXmckexTqVMnh
IlGIi42cBx3eg/k5YIn5rb7U3pb93bbb+wL1spqJ0AdDPpeGnC21t0YQOyzO2Vkqx2etNZZrtKAE
zVnMFydkzEdYS4amN+k5vm4v495jHDJoBLril2M51EOazMFxiy8CnjQwawV3b/Uk117TvwKd3zJZ
B4QCfwyP4Iojb8j+PcPShyP9ucfxihJVxaBkLiR2y57lrrAIb+endGmxulyhkvG3vH7LaNtx8CfS
yhnOhreNBLYnIhyUPRUkwD4PGg5+DEcMVNxky4nDgA7GF/6y82645+nctnslNpgnlYG5St96s4UK
hcQccQ85d0wGpOrLCBnDaHi5oCWan6batbWm1bWLxMLfkEIDaAdgxjs1IT/EdtsI4qRnnVWXHTGx
33H97dlHz+xRHxk+rDgABUUR/pk5MDzFnVQ34rUzuhVYofFqvA7YVpO2VjLezdbrxnZQPJ/rqRRp
Uv4qrsWlxiT2idLu1OyTiiIHiJ8YJaPL33TMB48zz4rD9Ulft8Bs7yszXwm+1E4OAppk/q8dRGh4
LQ9P2hLn73DHekm/gZx4UHRx4M4wmSiPtneWxGEQNK8nmxaW36TDDfz/UozADaH0QWtqhLoE1O8L
2d8m726T3tumTVpwLGxtnfNteEtcx8xyuGVShdy4C5nD9Vxhrcy+N5y+LXUCyAyKC3UZhMaX0nBQ
1OR9oZxxppI/Q6zBS/oPnin0HDRykoewiJKRTo7rswPJqVbPO7Fv1T0aWpYONSEDufYz6efRd5PU
t38xFFmOaQn31ycVWsaaXAIOATNWfiJaWcDkLNQdpI8setvpvJOivAD6f0VqXb2zO62uAhntkhFq
eE4NyYsS9d10kBHWAuQnWvG1TG47rqyawmjvrNVX8nwzKJuK0DIBJRJ+85LkKluePk1Y00DJDs+R
MmBPahh15Am5nfo3JgqYqcIi1vFrf1sgex+fyl18+qTNw8bDOsocSNA0cpkToM3uEbrojSF68ZAA
GjoMoAiG89YLD3N9kZE5Ag3Ak1UzF3LjpFfMGoB2g8DypJuSUwwOnCp8ksbD661rfD6QMb1khaSv
H0xKjzu9BkfYQ+N/TUitLx9UMmxDF+TtZIhvge2SMU4xQ3MMZsRcHpZdEG6sEHNYQok5J2Tr7GxN
aPHOQ5Q4OV2vxndoK9aNDa869BIFVLztY26fQ9fuejCB7OYxi5/5XPP/M0rGTtugkq/3gyxZb+XJ
Xvq/fiJs+iqZ/4Y+xpmJPLgD034babFuWUNrBypcSiJUWKE7Bzxj+kiSr8jMZjUxG27CFYriQtu6
soxxY/7OPvT/Jq4LuFLN3yngTQHlQXWL4H7Hh5JuuKj3kzXPtrwk0zmuzIZlLZIKharXXt7j2dJe
w4p+0aowzcKBMiDgb/BQIrXJgndfINtKoZl9XkIMfztM3r3FbJBooqqfz1ABktSonq/Yey3N6cq4
hizDTzEX2RqpGveSGQ1ndoiPpXrrt/6Eku5JeQJvP9y0oQ8zd4NZtlhPKUPkBNsO/QBTpomUBWox
IZNXaANrnqxNacc/WuGQf3nkOmh4itYYxoJSz6yJi6aqs4xl+O1/KQ+Gx0D/RrwC0rnd5eaMSO7h
hA5JXIK9HbgqDI/U6qDf+Y6c9R04si/p1i2s3Ztbm+GTYusbjTpzPOLot2K+kkvm844vCLsEw1hD
YTy6iZINJoxM6iRBn2zKv3myj8CsL4WttZfjGCmj3gXNGZdl8Jj3ysKyQqK2dsfdCbwf0jmcLGcN
SbOmNSqXJowL9KhygKzmlIsMAThKbNedCFORExtiTfXozBLMCR4d6FdOt4IIoDqOxDRsEtZtPTiz
Hjb10NRY7SV6UrTt9dVl/zcI14Mq1/SxLg8fz/mZqMOieh1g1eBt7F3MSj0ELa731cCFOhpVtoH2
EtKOD6rnl7AYIJAdwpytnO646Qa+FkshcPueYcpESll1mmxKPDmk+RmhzYtmqtmYqVZoAKH6Xn3J
3CTmFB47O6D/xUXGOI49AxXCffCEaKsTXCabhx3yNkWjAo4Oy7pPRCD6OwGsvff51mR9IMV3Sfe9
fxkDG/gvLMxeQbfzkB3Tdo8Emn4pgmHBFbdqNovLbfg8Qp+bhCCWGchwqtJ/4mAK3o+TwRL51Vdo
LD9OWtcox+ousGWfO8rKJN8+wn6af6TOuGs5RwgOm5467ueOwA5M0sqWmD/GbBrgF2/OfZHXDlNM
1ux29BP2Xbgi5l1MFx8biRSImufLMpBWErptjaFjmjq4PQJiKvqmrtiEaLI55yLt4uiucppvUim1
EznXnDUxWTqaD+JTNeRmk0mdeXtdPBYCaHmMsx9FOZtEXd+QEBU32iGvac+PaGTv9vtFlV5ar8tg
h4fUGeSlVMMqXQVmh2h201GZLIvW+RjgJx43Ef2RZmNeOFrhNLWgj3CzZgMkdBldfA8CtE9NgigY
/LXKPprfjduwqvM16ojbi0O2Va5QqOB5TfZKUZsES3/siytDinUeJIjQA59tgzLQuEUhlTh09sTF
i8iUWB6S8RLnyfIft9a+QenaPKvbUWbwRTPTAfK9G/gG8q7e70GEJIfE80CLVLh4x9SNiSBk002Y
uwu6hw2D58r87VobvQr8ijBh8pYtHzYVJsyQ+hmV5KlfKyuDUw03GO+ce/AaSEvX2a0SrPR2JhV8
x93zIEVIm+dBU1QlvHUamkpkKXT07z9xHtqC1OXf0iRr+Mh4IeQltobuzUJ0cDAVPVKOcXgftq30
80J86wLYgHHPgY0F5J4lzul2ypCdP0OaMcjQVcMAEeuJa4f3IZxOoW1pzn6RxA15nCb8byhcgwG3
qHAh1eMdBa1V2TODLhx/o/aCVXGxowk6K3B++a/qlBfymhxqe3qSAiP2yzOZK9edKqddIG8Z2B/J
t2kTcZXnhZVmhOpulna3SquhnLkBuCsI28a2CdOKKYRZxKSY1JMf9AEiW8WnSwRFrswJLZrnfpa1
F+qU09ufeYdVeKyziU31D2W5LUUh6kOa6xgha7G3xH9estNEkmN2OSsMn4X6B+Ae2H0vVWnX9138
vkccLCyDRzqnDtasb5L9d2DvUeWxB2w9VmlILCBS65OyX8Jylr85wEXex9AwjrQDWj5PTzx1mFvA
oOeFMc9oSRXvW8NWLgDouG2+wuVhIECRtDHrPkgL3gLbtGtaaU5OERwpLTvisZvlKGlOBkdo4yST
eW6l15wC+a45WMAO38yvR6157OuRDje2zerqp16vb1I5eeqF7/al5a73t6SS63cKOw05EucFJQvk
XNI2VOYU841ljOA4FtZhixNZbRGvLUjNRxz9FZVR1f2EC27+wG53796TiQe5LN0C5113TW96dhAm
ddrJpZ9dG2akQVQ2nBj8QVXiMpcNAamoxXqe1PvUMF7h0sLBP/sH5nFug2/4rXYePJiwreBGT+Qm
BWFNHJ5O3sH8jc8J9DAR0qCfUGodiszv7+A1KzR7AIwlzEOLAtjBMPeFFyQxQWise7y2mG1uHt4V
PbPxfqwdR8LOruSKCos7rsJHAYODu1N6ncMzcqwskHESwTZby3sq8wd5ukRsRtWO9Ne/g0tw74et
XAiA2Eh7Uc+qh/wMfZ+GPX5j82nAAlJP0RZOjux0HB2P3Z5VYO1L1/5uNmCsI0nwnFKg3KBkXz6V
3kszVVlto/oG1vZLg0c/uG6JYvL2/yEfZr7hsAIeCkiHKG8WFl1ypKhEMQiHN3e3nlFQnJOvPZrx
5iXzarq1nKrrXC7HaJHn1ZD5+KKNqxGcR0jp+S34ZLUpczy41tU0RBYOubEypMu1FS4QPv/+WvG8
sj2YqHOxcpztNMMG7DdccKPj0xp/d7DNBrkTHpJIWXxY+NEQ16mpsFxkhXB3/OvwwUcHAwxY14On
vrDgYZSR1QAM6lamYY51Rp0lWdV8z/LSxe3XMHB5XXRdVh9yHM3pYnogeAnb7quBtJxKD5+YnHkq
qKIS6EfLZkxIlTi69sR3vbv54EDh65MEs+zTo2uvDyZf765g+sVVj9qgBE4ugyR/6hFy13CXdJy8
8WkLFoJ6OL3HW7AnFggimSdp057pDoeW5np6W+9/8DjT4Af41+icORL2MwjtNZGQZTAlVsCsZMy2
PPc3toWLCNGHRRNU6o/CsLsyJv7CyIDVS0wnhgCcZ2won6W9X2SKNE1gcfD1OW2nszxozj0Ph2u9
NKxN1X4sqg9HZjfd6xjeFP20o8LsJw6ZfrN0hGY7QSBnPddToLDkYAYgCsEbz9fxjsvylN7/7E/r
i3EZcVcUaw1WysrRVYj6JUh4Rfsf633E3jmqLpa078oL5mNH1mZp6GAifR9zrS7rDRzFncVSmoHQ
u7zuTqTuZ0CpJMaWayY5174htFczWno6lDAy9JtS1ZTQd23X2Ew2IJShMnL5KxAMwBQ1pAelnf65
h4r0mSuv5g7xlhjDZ1zKgOOXwsf5UxSmlGK32Iba3yJNvaN99+4YY3D4Y8rlC6IuxE981j3stRFC
PK4iuZv4APTYzHzN1zkRR1nwFTnOFrkPNV+57DfHQHngUHY2Iy7juB7E3dhPoalgNcUljOWVIJMp
zSvHk8iVVnSok5KAjL80wd5ZmLmyvZbrgx86vE7TtzINeirPaS0MwUkIfCVHtGmVL31FYAZSWZtw
ke7epxe9or6soO3q0nXuqxNeL9wuoK0QRQlDj9TZtyrqYtEp27j8SKp0OgDeltvsggOpAXa2odPh
nasuA+S3V3VyWHgS86mGt3Y9UNYB1IQD6gsGsAHnO6ANmBWNkUz1AKMEsEjYoVb50OChQoWCAjVL
r8wEIT4B31UHm+c7RuZlY0i25FfLCME6aBMMWaEXdJaqCn7vyps6gOyBpP+RuBGZlb67w7XtbC8n
44H5d7AKQHOaZMLc0zrP8Ye+sS8BbImHsDgPb0ddnpVE+IMfi4wzdissuZmHzWgDTBBBr6ZYhHLm
8QZ/1acTr+aqbhdXB2YVsBAJdJsvDijAsK8HTLjLNH9k5eoKtJcaLNUnLXKkl7LizPP7G1oZRlbI
MsgboGT2Wqm35/f8COVpkf7mo2r4lO2KUTFOfwvnz3Y0jT3ShOsXJ9WglFGoWr/2aaEcUtpxj00U
371LPDMo/kG1mpXZWg469Twic+0JVpayhkODtxrqUjdvhKyiJhK2q16BeAuePdoTRnMRMVttzI9V
++p8bbmNJaEZWGDD9C404fcPkisEyNZywa4eLGpNRo/x3In1EJ2ydxgIlxdHoxVaK1aPJeORscMg
T6WRdjpyREeiF1kGxSF4zcJG+X1DkCD7FPQ2Zr5mlwuG69c+86p2fFcg6TfU3mZPM1mlwTBddE//
E2mXos9jR4wVAbbnno4TGeS+x6MAM+YwFynW3aL8p7WOYinW7m9LQFtCeJhag/QAdHRmRXx/ipCx
pFzfTVdMGysImP8Mhv6asHWM6dEOn0NQAkMk01GoZbONn3hg78j7UHVRSzNGh1CxFtMlzzJs9B0I
X6L/iKX6Vd+D74lMxdK0TZjqkZawof5bssaF9J88JKUIN3w1rDXxdCz9D1eVhOvg/kIiacozC9FJ
M2joKt32/Rx3nBhoTCOQKSWUwhEzniH+j98Qp9ihCkUseGkeZX8N+wtsfdxkuUYcK2bhqlAJssBv
v3Q2kMXU2po6KB6oNEH/4JRWQvWTJEl3eleRDzSBgTC7jQWUEvzFYeIsD/yNZ1yjg/EYYgNSbOBw
zr2vr1MTiZoIslEAJBxQWjFmJ7Ba7mO9DXNmgPrp4akkZFOZHKXkF/bsoozFfuAoL+Zgx27aKn5i
BZG6SYs1FG7xBjPgpb0kTP2tcXS+TaYSPoa01VHtpZ2jQksI582vuiOhdKPgZWM9Z3XRqepeEOq9
SIsUZnwPLAOjsIZS8HvWOrT+ic1ry0Lm/nRfAK/Rtf4/zCXDoRloYm116lXga+JRr5JSKO682s6y
AHIPPXARcJ4NSqUgrV5V1viD9gnLjbYPGxWIMfjkl5+xyXyGMWWBTUvGLK6Fak3HluYGych/D8rR
hrlFydkab920yTflxfdYK4fYwdtvx5Me3YeS5XA8q6dUTgOHvjBImlf+K/S6lb5DZTkIacLsP7++
xbrzcMp2AoHPuyHL2Wt/5pOVHY8CIlw2XIIW8Y44YW4z5B9CLigEFFE3opOkFznYcJ/0ZmVsR6f0
BsI0JIv5bLvh2994rp24W5RH9EDZApAmp775A3rwssgC63sTMLWcPCtdNwbz4vpjVhADOkOrD28F
AHapUN9XEBCW+kEcMCN4Jfc4y9hh4KADyJItVdLUwGRzO2rJ/wbX9tKV7h59JIt9cRcc/K55MKAo
kdPtyk64U8mkAbYZSwKaLPw3aLNSFIsiPflfcFlUqF97OFtX3/MYOggTRY+JVT8kLYkIH/1RvOX/
lb8ZZOO0t867Kf88Qx8crQFiQG08fdD9heu8M3YbKN8Cw0GmBp8tCEto7u5IYXL3C7BOpXqnyicw
YCEc6MmMd8pvaF3RmIQHSVA3xRK3dTkbOyU707OqdRzAoshsMLMJRxKCBls/Yt6OUeGHiagYlwZC
gF8RKsrhFZIxfiLRaJ3IDHn/k8EHTrC8q/Co7Eb0IaeKRw9DD6c/qbkJLwZXnyOeOP2FpGkpbyuW
I3rOnV0zXSeTD6x5NfFDj1aYI4TH1P6gKFHWAqxJIQbEGCy/8vEKwOAQzl2wrsMz3AKX31J8QcNy
5uRHB7lq/7OKEsAYXCRK3YVqv7zJe4ozNUAtH7hQSKisk1QoRCEo9SCwVsIqFto1mzuGbwp/5lIB
lW1ls6kfDptUsJqZ5cLiHBAmv/UD+iUqiLnHMfBI762aRt12UZGN51yXlFCt2d6PZ0HJfn+cGDN9
nR9Q2CIVQH6yZf/1ue4mOK1TvbPCatXj1VhC1IgEGAS3un7Cp3sIFoBdareczuJJ3SALeavH8bz8
BxTAyrKa66/u2J/q4S0qfeTVya+gTOXXwaMVymSFrKWmGowIf6DQQqvOyYmEGrsJ6vgtrKkl5PnV
0BnquI3wfHrR9iRrdRuEHeGTRAaOnvpAPwEDSqFyJN80dCdhIWKS5r52S8Yn7J6uPVYmcCgXnecT
vkWPGBNDY34HVa4dvnyYkHdijDmP5QQoJ2AJ6oIuReuUnP5PzUejqW0j1wUcYQw3S7+CQQh1PKvl
vR0MQW8nd6Z+m6aplzDQMXnAzq7sGyLs3dvxyb4fZiphR4WnDDOwdPEC06CiTdKI2q1Gj74+/Jh8
viAmntOGwIzDikvpkxVJlYYOMsQLFqKjNPWQLy3jdkeIqkPieOu7CjwirpOVytCI7tdOtqOSvvj8
BaeujGKnds6Y7wJ4qYubj5cGfg2m10ovXk3v4Yerjhl46SDG3iwLjwlJ3o4vogBRoRBiyR6iRtFP
dYcRjJqoy0WLbWhL2e2kjQAUdnXv+rSArvveL7UNtDueG2+dPnUsmC+CsF/jz7gZPbGxKX1JLbmD
/cAR+AJxrfUM/7CWDGTpRL3ekUOUSlCmCdTNzXSe2gjDkAZQve2QN/qv7c6JmcYE23NWzJ3znVxs
Eq97apdtCN6HSJmrxP9AjzZBdgLRrgKjq6CyR5JpA9ZTwZuvGm1cnWN6IpyJMfrwVKMaW1K9bQoh
BOeFBgcjCBL6v/B8TBlAdChFNWkZhlxIWhPgu2wwKRHGi7h3kvDO6HAVCo2zLi/eEWlgoD0PGBm1
TV4AI4TeeVB8byGE/GtJJxAMqQ6ZodGxwEYPCHQCk0Tl2OaRNlKJRhT5J2iQhFkRqBIMxqzBiTPI
0p0edVb5WgI47oT7DBIQY9xB2M5/jLYRGPsHFvSemXHY5l87GRIsN4IgjCIIN5+Qi0g1wgXkhyxA
HX0goFKlggB3/my55kE7nuRxDRNMttHM2Bv0eT4NXZH9xnu1vOHKFMXkGwSDVj2CEI998BABukdf
jdwjgY4trmWjM2P0VSt1H28hm/FvBioVHbqnrnhuigCXROb0wtpJGiBENbpM6/xprs6MK2bfuIKC
AzaW9hG9imV0TEEY3VpQF5a3DpqI7K9BHWrPBs+Mllq8CwkOd66GP0OC6mMv7wAVthCfENyrH/ar
Nl4CDHpyelhK3k6eU0/xB88d8eo69sp2aEs6MK0onRdu0ooiKpDY5y9qbwbzQs0q7cl4PWBeUwTg
kmsvnYzRR6QlIZ1iZPC4tkvLOR+BsqQXWy0IRDS+0JbJX/+/w82lgAqaIeHA6mlBWKxLotIoBPgv
hvrju7y99zGHsyN2W86Qx+6HawNnyCUhyDoHz+tWh9q0F6+Y0mgWCk66jqPMjvxgf9kn3rsO7Do2
NyKVeh2X91rso5LzMdW5hqlUWGD+IzkRpH38j19aRgIlUKFq3NFhAPcWOLFHeLNzVJYGJRqkh47l
JaDl04NVSkXv+6GnIZTcwUQjLwj3NzSisxcQX3tq7Df/yUn9l1CuhZw0x7eO/tmyBT3lkhGLD5wv
9eyc0laafag86aZXT63qcz3GKSBF/jQxKf3PsUfGqERgVfHnukWIwZS4lkC6slYsvh0uINWTogAW
lcXN/nkKDexscJoeBueduPUuAggIyFyXGejC9E0ZBa5l7OGh2LcTvEl3AcpABDcV7SjFvYdGqWPa
KLsCTrFdAnWJGkLbB1xeaRme7l6hy2dSNqjkP12+tf98tfNWrEV5Xi5lUrHy2LF+ZWed41nKSIw5
akdK2HeCv7uyshOA0bwxuVVTr6YRHGRKGAh5Ifi/zYKH9yPRWud1CAqNHHUOOiAy78jR4k2K2tx7
B2qYLry1WqGVs091mpmkvNz7I+Qjz5s1JtdgYGKV8zCq2cNvzAxU+tzoEWw+1ckSOLtI+kQyyWNq
R8TZmnZfRf3Yq5dHk+svh2AyKHy/P8pfHlj4o59PaZr0w1z7F0M5fW+C+OrhAy011n7/G/GnG+PL
kXvfIQSsfMN+zr4HELehB12GC5LxMRkL8TY5NehGqMfeCtm1Cs7O86ZPO/SILTTOJYsriaQHuyqJ
OaekxErL6KVJAEt6CqxXue9JBRoi7JJJ0JwQ7+T4xydzUnopCOBed4VWDr7IDTEvsY38TISUR7DD
5kV/asphYLp4FmhTdep1lZ/1d+kDN1BN4EPMtPzUSdtyOvTXTzFvIS1+jK/Xg+kCxevdrq8C/3PL
MfF96dX7hnUyBC2H9tSGRy4yYTHNY6rSkOIUkscgFeYYLaXesZ0nqogJgKO71dd7TplnWA5+n44z
tq6ErqExy9JmbHmmkMmOsTevGrYWTkHk2HWWDiem5GJblIWj4TbmslMZcgtud+2liHj8Y5J+RYKN
FJRlW+z46SDV7qWQx+CQXhdEIFdh6Bw7RvaTZoxf/Og2cvRL1jK9ZRN43qmmWVXgxqz8xkr8HXRJ
vfRjDUdsWY3/Zv937gSJhRBgJKL7wiADTeTka8an1hM2hRcvG4pt3a1hh7VNxhdc2OV2fKEkUQUL
aqOVeGqXyZpdG1t4PRQEYZvEzX0QAVIYErptC4uPS0RCZMIyoduDFDBf2yZv53VdtEBcy9fXx0O7
rUGV33IlpjJRFqi8PiUtYblYDcF/kFkDC/PMh9ma67TYzUTVz9omBW0ieIYjRL9tYxHcWkp1+ke6
d0l2zets6TA+ZxRL5Tc8RbGOmiYyT0YI4O56MLFSXkK3nIK7aYOg+AhzQiI9i4vcJs4DoXc/2yFm
MvM4CxIDar7xLEugYjCW7MPK92biG0GcrnX7Mpk6g7sqv2YkbcKN41h1lWq2kTkEnhDrtkQnodPS
ukBKJMBjmSf9o/BVhP8zoxKcHrX+MKkjxSGgbuLS+HkYFSsxtVtZODIah3SED/46TugBQZIALY0j
iyuTHmGzI0HRwUmvE5s8GWbl19KJ+xKHo8pAgmhANesa18J8ZjRPJgflAPjOjumxX2la4RhEgAB8
BeUIbid0fPj9IuE8xoMTW+vun2y81ZiqL+7bPxGqS5xs8qyt3taBgQIb/v8I4DwVvKTYKj0fk9bY
uGMdlJoPiuIPZ9PdQW5YzEcsDoR5wCJwWIaFxYMAXWBrQxgmoWFs7LWcgxnaXh1Gfw+urxSSe9B2
VdyBQcaLoCqueHR4q0MbEM0dFn5dR11bJBL+7fN9k9kdyJoxXly5XDk+y0/Pn9rUqfs7ieCOwJXK
ALff76KS55SUJV6iQ5AqvbQfDWCWx226X/d4qhHGy2lvGYD+X3j+VC8sg6XpARbiojziQpxsbvxz
QKIyz4RGT6D4xr/1IWb5glhdXsI7mR6Hoon/eiMt1oli5DixAIBoZ+v2hSTgQ/86rxFq77ANyUPt
M4sxbMkiF9yioh6cyKbokKKbt+XaQpekRSV7X1ifJ7gQ64SxkhaL9dR0Qs06B6jIFPKEKarMsVJi
u3dSrmuQ2uTnb2pSFB4B9c3s8ZkRERlO66yJlgfvWyE9KRd/363YHHPyOynmIOjh3dWafij5ZF3H
tNOiwL4QsPLl/QH+7OfJMip0wM+yfqMjAHI3mcwt4awPzAINxshekE5ov44fMZFG/iDB6R80xBYV
qwMatgQDGvcUPOlHwucDoiDnSop3lc+LBj29sYzXkRHoLdqO/tEqP4Vi2RFTd3MuI5whSJchAZDn
LipoTUr5FDLsTn5Mq0ZxGi9taydA1omBWLRRr+7tZTF/c7XwhHDyiAGFVJAJ7KwqRa1N5mfhls3D
PERJ5cM5bLs98LADj16D9Y6kR8NHORPsXXdHTz1Qy7+rCeKdvNpzQK1U0LMAx5aIEKKvdjQ+GGoY
NaYetkjR6vdxYHWaIY/qB35ki0r7DQ/zvIoNA0PPitj1Gu5kZ89yUeb7MhruMVT0OtUvsLwOCrJX
P8crazvnNAVRJC1QzkRHd25S2+/XcjHa4nPBjyxXnvsTaSAKXdUUBQoQLA7wkRvird2vgK9G6nK7
l4SMkA1Dr1Sy0v2sGoZZNJ7lYcTKdeMecihQ/ouUJ6E/i5Xcc7XAMcLcYaTD0J2bXoX0yiLAbciG
4PY7SVq8eu2dWghlYnvV7QaIqWeMT7YLGB47Dx23jnksGJimtED0dr1IETpmvQhmbZ452b2838So
7+zYTSHlw/uJXXEV+qrIi6orSNLuCCNhYoU7+mn7GySvdV6DG9ScqMhx2p2Wjik1FLkmbZ1rRM1i
lqo2bc596geXVmhv8h8G19iLImJ60iiGwp3Agg4poYvVZ8iqgLSz3KaA4qmABJ0kIptlcHURg0Ug
a6dl6717SpsxnUiP0ojB11c9gtoXe93e8A+b2aPlR9ylTwq+cRiHI9VmeIvdeXRi0FXCxhzeCoBM
YmRL1bZ8MkdovV4cn4xlUi3Xv76ZdsdwIaoQEQL7XdywARC1oYWsDmCQi/6vT01XoFPXwCgvmj6e
U31Gco9Kt4EcUL/P1XylA+Pj/+DNSLIAkteNrPp+mjbUc6HfuUBxo6RL++QeGzCmNBxHILeuFhs4
l2LEYz+FKZULhU7ibxC9/DbNLyY6ulCQFx9tIuZI5rZC2w5+foyuixMUk8XrmS0PHjWUtfWgwBYh
mUHnq7I+GOlfQwwBzWdkEt7c1KlBfc5wO21PaKNfQHgcFgxFtnOq+dbyQjQ4Qdf6Znjowji7cpcH
ZyAXU20oOt0A+0nLiVRbSTsPjHGu1OQnCHU7QiiYHMH7tYBjsKZa6Xz8ybg12gPxHYZOAxCrgHwG
fmYfG4qMmACSFQLKTNrfQ0GviSug8GTvGINnpr/RoDz58jAP2Z6hEbkGPaMlIMJ4rJQd+JGB+2AY
kB1Q5tWNt/Tp5KaGgiu6IlFVlg1nSgPqlrPNJ2dihimA0cG2UPrO4mHwEByHVB0AEQGsI36t5aSt
wABE0Ph62gmYYR7lY5jHHVALUvN+tYH65Tanr6wNMq2cnuvK8lbLhuQSCop3Hhjk3c8pesOiHkae
0Ua6xtn9NSxQx86mB05LcLQf9X6FPX97MHfghTo+rKchLoUDdlZK0Ejbpsb34mT0wvucyOpkbnTK
pqoXDNWezsvMbXSgMe8UZONS6nwc4n+Jge42j6UkAqgvDK8VsmlEkfEnvscPsJ7gJKaRivGuuvA6
mGIqbf74MFxJfgXbjN5lroO4OBfLsp/KQ/2vfN/zyZltdiSlCT9RGTsHfhFe7AYpPDUVV10Gojk2
NNS+ZZpqc/YTUQwSzTdCRc/7Le4Iba59An09sFfgqln7jWaHuGV0+v9l+cs9k6a0K5B25Iz7zWAY
NJLmHzASXSUiwuVQkIsgxvofJT2SpKsWUCvjAZGapJ99vz86amXqW6fjFwEb0ZcchVcVt3wlV8gE
Qr23PdFYMyK8rOIKng/PHjeaSkdDy+Q5G/LmnsWafrxM7TJ5mjZaR7cb0TMujWYgh+klYehbaFbE
WgyU4kUEYBezhjQEXB70euGjEvpv7Ak3M1TQoKh721dL3X1Djzh8kwOgRmp6g1MKnF5BuM6DQDpa
NMF43bwgRHE8v28R7IHiqNSVmeDoBXd2EowdbIJxc85pXHqY1Lge7tIyEMFUexjuR2Eg+6F7UYiS
WDO4ELGqRt0X5DWadsNONWGBH2kc/yCMCtkjDofMGyd3fdGeku61HI4wD3VZ60J/UBK/UiyGwzxF
ZUjQZuf1Foblq67APCldqr7cIg2SBpTke2m5ZQ6v8NntP4k5k9R+0bSHg90lb/CDyap/yalBGgzd
y1AHc6P3PF6eWHHe6tAI7KJrb8UO1XPuoJh3bvzGYxA4+tubCeQX7xlNBLeI73ClYqJ472hxw4sF
Pn0SvicvnwIFlV0wRvZ1UgxKEKadufJuBPECtLZwnbCqxgJsreU3PvkJaFFcCoH2e2Cz3Hsjr/kr
UBTaBv4XmnoEl6UwybvxFHkFt2fijAS4UeM22iGMCCPOXj/76N6xW51XIBwJmZsn1SVcxdblAfkk
RwqVH0jIaDKz28f61IikbYLZ+AW4vnZbqSFrcjcyJtKsTrxhsM7DcmbWA8B7MR9mqj8auICb+n5Y
bL2qnrjO50pkma9SOY3tmN5+CvpHCkM8vAAka7S0WEFxCx5jUFlYLQDxvFofSLHzhiwnOEpJ0CM0
VD2OUFhkfjtyy/0N+5WhnjvkwUzJMH7QA3g7bBpqGPnW4cbGn2+gTI1oQxUbOT1y6JxmUZnG9NMp
DVQQnOhZS8lzezxdfwPkVoPUeTPyNuOYvpRTpUEtQGChNrHYFcYmCbrKz6QszokZP41Cj0FKZFOA
fh8kOJEA4+rpd490c7/yb7pIOkvtqDey+HYtNSxWJWVqvKbUZGq36grGH8qtRbwaKZPWpBmvYx7J
IORFWZQdKCJPQ5W+O+oSpxv2DhazxWsq6gCgPmt3JJiXjpfVEFuHYf1F/SmFZuU+qikj2Vqyswwy
6cyeIT8aGOh/GzLjUCrB7pwqmufWUue0bDMDWkt0pj2QpNK9Kr9om3FdNrq4c2UuPH0oCT5auHFP
xlUj8z7WjhScYGkQmw5FvTSHly64xkKCKTL3mv5hyzG0rIPS02zvIXskpVCIzZg2ChBXuIlvhjUA
Wvqf8QYXtlSELiyI+3ZcNpxt3/ipFii87u6Xg+zvO3TFkLQiIJkqFRZKz/+WgPTq8ckckNahqVqT
FGBmAWdDuxJCsu3TrpSXl0FX0iXtIneJQR0Sd8uWEb3HBXC9zeEaSb7NL8s4Diuveele942DS/ht
mRvB+522Ey/sI/IRlSCjSOFiGaEqnwDznF3zHCCRSrkbu2sX2QlkNZSIhBltG0hA+UA0kJBL3HAG
ydsK9xPVteGqtNcYhNzImU+yii5DLIu63FaQDr1WxqxTftFxoAM+XSdBCaVpKYgFFS+SuIodgVAI
1JwDhoxG9MTRRN2LVcZDT4VRymsJ3+xz3wISHxVX4tjd+LpLJelFPAP/LwcYzifG9gUH8ECtecLP
j6leYnqPOusaNzLcIx0BjCm6OQgUNZnIEtXNI4OTgZaI1YfccyoOGu0u8VqKzaI/9aWRj5rW5OUE
u5DtXa3bETLacamvX9eiZ1up6LSf/nhCdMbHjmEujOPkoxYi6/gwk6gGkIF2xvOOCjjo4VcFyhdZ
LpbTZE8IJ7v4AZLYhq3mQb048qZSkQs2YSLUpwMshOjIkj1Jg/wj0L3TmJ6vV8RTL6W2Y++F7qfD
wX8dKIcGzVnACl4nYBIQS4i6R7DJtZ/V+LKD14dQ+41lCWBLZAZhZj3LxeubhpfJ/OBc7QvVJYNF
k5mkf/i7Zuk25YlVkM5qAShCMyJqlqBdYe4ot0JPtsd+wXhKrYD8oizjQDNMNgXUcRKbMCxS3vU6
elL0Ig71JozXAUMGqMqsYgTIR1k/M+rsOJuGVLjTszknpiGzKCh7bdDK2/f6pavP+KJ3/s2Jl9S2
OwPYnjDMf/ce+OkNmTf1gZOeTSaTVlXm5x70+eKBTOv4r5o+5x6ovbqJhXM5VCn1WI9ZNnJmtOmK
iZl4//vWLpH5QiPoGicPULp27kjnV2R0Kqr02m28kAi8O655NPdzRzIEgjepJwhVPE6eQS9uglZx
c7zdgeyarY+aecRMxqVtHZUK3TnnODzK1NHRUImFUHt9r0Rpi1Q5MvaiEwNbPLXsQrgFPMPaX5eL
C4whrpGb5dxFgCBFQ/uZUtUC3k/BZY1xQ/aZNIgriErjHx7xpfcqkkF9Dw9VkNi15KnLSM95fRfj
OO/pvAqi4t4laKxweh6+1T0suj+ckcbdoOIV90Bo7TOmwwYCxGeZOZBsTO8FddC68dcGHshc0Nse
CsQfX/X+DeA8ppSE35S8z3u59lrg9SUc3YeTi1Nr/vnwmKpATvSqHz7/OnXTAN7jwl8oi5WeI9/C
lYtNyAl+424BnLcZHH8cg7/L6fhaoZx12U8JdBfy+HMm9Mgr5BF5Wx0ZY6ijhl54+NBmtuQokc/v
k7RFg9jb8eaw72ZVpQbCxdhWR/yGeiG+1DgzucizrjvvWFGK4d/7nH2IQ1iCCqNgQODVQTnjYLIs
eFP8rSa9pzQmhYSPYsAqz31fW9BfSi6jFgit90PqCZ4xNJBJ26BFZmO2aCvztQEIf4AaHdLoZU3z
XCJj2OTreLTPclMmSBuxv4+HL3EkB64cqVS8oXMNBzNLYVjnsMy8XDVo5h0O7DOdQ3SE7S+C/Fuv
fXx3auqaBWgZlRGDyuUIw+TzLPdQse1iTBbyDq9apNGdVFhrKb2p14ljpx24d7ESIbnAfcuvwUkW
c/YuGIl7wh+ly6TCgcR2vfHq4BIe01C9c4ETz2V6b5EOQ/CKqjTfpBkUXL73CnMLN62bkukf6rqy
5EqcEcqZaarrJ00V+G+hr7+yOyawB7XHlZDlK6Gb8i7jUM1bt39WWn/uOAlspn7pJvqeasasyzeO
VphD0eNPaTboVAPncjUw8tyJyfcEbZe4QV1+fJXN6bwfkPmmAwMJAGtbLfu8nBax4cmnjskUoIA8
zL96HDcZgP5bn4giTTjz1371EM15dN0cg4POXgUJ/zgIHSd3ofgoZF0NO8zZWU6ARQHc2bWK3jf0
M+TYeZTmB/diX1o024m3EzFlvmcSx3glDjrJMng++iA1RW/7WwcRxi1fB2GU27YXCvwiSMLdOzB6
ZTb8z9FCjB1LXB9yeLuYhDFKYhumCsX+o3Q7PZJuAc7Ckf7ErNKftjfs1Dplzf/LdU4dswPNjHov
M+VK8O4T3mOCOVEONddbPDKH7VLsmfxY36y+aManGUU1fRmtzdH5uDmZeChfQuLZ/4Bx19Nopc2o
YNYVwzKRFs2KT0lzjFl0L5PN874ug37MW1tTVhmDnQQLRxx5sK40qnee4Fq9HL0SRaD6Xwz9KctY
/EhffTY/MdPkKgU+5Z9EKJ5WG46IrQVJ81yycsLbu/vUiES4gO/x5dU3UEh7W591EFhzDmWXQbeq
Cpzi+tpBM94Ir6jndZ+WqaDheEHfWs3ed4zWJWQibv2H1oXEk5oQHvSvQSsPThmmKS0Hw7mXoxXy
hwo7oT3MOKoNvjj+tkx894O5hnI6u136rpmPmE945i68AMsxTCLVDkWR9Ca7JyTsSzT0Ndmi6lY8
keay1bb5YgHK81Vg7jqm6ErVoS4jcz6ORwqWDKg9EELxTAITtV/gTmPslsCFt9b1ykctScg4JHIF
n1kIT4/n4/WDgeuL2TQUSxwl10LnC65vAkQ4htEIGmcg470hk3XyyEP76XZ9xO7WChfEwcR6xypm
WrgHZEtsI6MbUPYehfhB49n0Ch/Pg59283/b9tg8BibYm7HcaBO07OSvO1eOxURbhMe2m577iCFP
ZUTOhC7NMpojJBdhdCW6P/yIaueHWliBCZLSFQBf8Tty0wuL7egi45XirnWuyLyyQAvNU8sqwrmj
7/oQ+bbvLZYakZE9qexCd6FmeEJLtpGap5Cm9jCy2gXU2LZGkEczU/FaY/Yk+Ol1tWznpdk1qkS8
dusoh/Q3qiPItg9p+eFMhrrQXxfN4Zf14M6UEdLPlg7hT2g03pqJiDWeZMMH5QY9idGWDUcLX/fz
z90PirPxRpriwS+DxcMGbqomGfY49IwxZoLTWJOzKQfgBpgeZYM7LSszsf5LLODaQOt5FywxYgU1
z8jvCWxtXd1qf44VJiqOuGglGX/mwr2gxd/UNbQpcL6B74avj/FPjpQCWCdgsgXCB0upyYP1HtZy
1OCOxR+jq3rp3JKZW4qaMWlMsBmpjbU7rNKcLhwwM8U40pawbIbxRwqUNgoptjSpvYRK9iHVR619
XC/0y0acWdinqiSGVYOWvtNJhHnDlYbbVRd7/WmO2HJ6fiv0NVunxMxslk5OyjLYx2dbqzSC8Dvl
lqKC4xtvOWCSCf6hVQ6Hqwb4mj/+/Dmp2X8S/g0c3TQ4Nz96EuGoulKvEc4rwbwJwIuQxvptzOjU
7IRks1nisgC2w88Ym+x7QJaAsNe1mZD5oATaIUcfov/h/jnjZVmkvf6gUEYI/OmpniNOqCja3Fz8
rVHzXH7+BH7EGtTCFC7eHn1u7qbfAzuZu2zd5sQ56iOitun1Aj7795/VhA8Omybxdh5aibDBNgBG
/6Be5Nt8hfykMZ8dFMA4EJfL/zz0Xub02xyPwtg5exOo+XP2rKl/kIifdxMo0RMnEI2tr7n30Gne
R2a0JQheyrUJ73AlQjoQ15I2FINtHjmx2BxWCNc6TBQZzaG91FKcf4KdRflR+t2plHAZzbwh2AKC
DV1gx+DcSp7G6F2k2KOK7UFhqvIX5sgeubw36GaqC7cWY5qGn20tKYTQSGDE7WFDHFlPfFfxs51K
MuTvWSCGOetu55x2dOgZewWRUerMZrXZa4NCt0wA4D60gFDalsGmFTTqWCBbvxeodNONo5pbsZ8p
5V5dkyUImDdHa+Qt7X1TuwyWD1PcmcsJOOl4rb4mChswatzKtBTu6tkY8YQuo6mHDWugzlA+RsA3
L3AZethPBR7KjEQgNG6nTJRPJBXQoyhhF05fnvHjN2dfsfUHqnFDzELyPXXhzkkcJKjuE0Qfx8LH
Kdl40AyFQ+e1BSuundbzhIQ9kzxO4uwuHRmNHGonKaVt+793DPXG8HKBryThpPZjahwcanXmLEDb
iEfJvUCe0tNe/8QNI2ME9YPqvFabGiYlnylQBooHWXgDq92t48rcYb0euoqGF4vQZQKwnCM4CCzz
Gd8W/DHJ7vS1qBE0zyMTbW9pncAHC+9/8EGxhk54w5io1jKeeErMMfPD1ADKuyC5Vdcu2ISj/WUl
qyMfRic1TN6a9qv3J88dwVh8aCICxKZvgVYNerTX6vcWL/lggSfV+C/lyFEEwFuZIl/Ucqou+G1W
Ix4dxsascHi1g5BEOkBHoZdligWmMSxTwJcwlN57j5ipxqx8Wf43lM++zGt37Bt3t9UgJvcsaBUC
MYjl3s5q/Q7zVvjDjuej9OgZzJMOX73LR/97XsiZVcDYi7T9NqZ1xbbooUvN3JB5ZnkRtBw5RzCx
tdpb1zTc0xIWCYnEAb7te5FopP1aPgG9ukBqH5A9J+4eDjQ4D1YOi6E6474FRc5ICoVRyZ/w+ar/
YJnsUAR+hHb93HyQBplbOW2gybYrZsxhkByvuckwpk/Y9uJb2m5ddkYKNmvFxSDmGuNUp4x2bo/H
f3P9Cu2Gmp8OhG77RRELIxu8O9ups3LG13SQZSufJSoULyeyud28TesJw143wtPdgugZc9IbCKss
3c8/2FMS5fUGbX2gaPI1Y93vpsYtSDpCVWP4x2slDNeW5QDMFJ9pWcvJ8s6ZCT99vtp4/LP0NvvK
oRDktssSaukT/AuVnXQ6XUcbpbeETjOGLdOR3yj6v7cncTgw0fDBqn2OykWGVSJ4rF9GurMiqJdT
Y2zMBkMGWM42SsR6BtoS8SHnZK8vh3cm/vt2sFZ4SiB1YMQJg4mRbTUvyY1bnIlSvteLihCeobbA
1iE5406nkV8Rb0diJs3lzYj4yp+dAtaSX6OXhgsPicWdf8SkVwb/ZgqgzbySrm4KhYp1zh5KOo9g
SZlM4MZfPKKhOd56UoZW6MHzlOPLuH73vkGKQ9RpE2BT1mKftNFFZKEuADE92zrZ3YodjhZrzHcF
iU4O93puXgg7vtsFdwIcWgAWwPHpl4ZvMljE7G1WDSzdm4+7BbMlvgrKiMCToKWg8gS3KOKTWQSd
lpEryXaQI5s8kSgundbt3TgluHbR7tVyG/qCtYpAU65+Lez/PtkKFpyTP5QXXDbHG2DqdkS3lTws
3vDwidDuzGe4OUUFXyIHy21A9WPCcVqnQCw3PIHf7J4XJ89XLU68FymVOMU17ppO4mQhKKNLo0hl
LMW9pUHnKpDirPP8z6IdBjw2o4L5XeCzA8baWSWFMdrPJ72icUGUTTj8E68lWyflScrxEFvHSiGo
BWRWxXl2+DFuxvGaETEpbJwYyhE1TLeMdfCFsNrhu0pI79yH7G+wjMXvF2vooKgv01sdhmqO62KR
7P+2sGxMKsZcJ7Gnx7VVmN/0I3HfJlV1YZa+knNFOgJkAGOWnWYp6MAE+iQITW5sZEHR3xrZTC2i
bNzw2CcLFsHGd73Y6HYWBNBVJmpHh+OGq6v75Zh0ItyeUH6/8x2QV/M0sce0Q1wiNFVQePORgJrt
0vJcV2cQyQ+3ON/1Ty3JiFxEG+Tv4grbJgojRAxyu1/bQwYFR1tkfXkbgo4/T2kC6fTg7PuwJnXt
51X/kxMoBZKr8EQiwRHvnuiXsIDWW6kAHQxqymXikQgH9fVIkoFNf19y3+LyRq+kxIxJzU7LBPzv
VF9ewmLKPBI9h5RyyhoHX4yipIwUQ1fsX/0bznlAsDjqZtpHQOrS2+cs4fWfkApcAR1kr8NxcIRi
pVJ9KWYMrIuwXezApKnHG+NzxlWzi3iduMzx7j+jW12jQNEqkyB7FR80asKSHeykTecZHD4W6YKX
59Sse/Ueloflc4xm2YvWt5NWynfstUUj/6f9WPrc/fMS71uL67/7BiUSHkxa+xaoMOQyGM+EX5dV
6bTIf3ZWVNTQprTutoIYtc+WeUS7F07HbedxQtURTOyJnBku+274jQft1IVv6bPUQmr64Se0MwUI
hIl79R6ErML0KispNDxCaZrhX3EsRs+n+beW4FARr0x9r/CLpVtBw4SIhdIKZazk21FwSsTIYU5s
2MxPy/rEHcm8CJRKT6eHLR5Arcwf8TTE5E+bqFLxFm9ykPFeGfbOr2QxrYmDU2IM/5/aHRtCqkT0
KC2QnD0pzbsE/vBiBfw+VDFkwIhi1B7LPeKzpPTMrd2ASI2S98ntcO8D17EvyT+mSqjy3k6SJKJd
a3narweMigIxFhjvWwvzHWcQQfwCN+9+ggrrPkKdkapUlnFDXatIIXHHvljm56gHr9FLL1cyXs+7
nmBHOzCpaj4F0CsW5KkCNAQACEJcA2kgmzU6LujE8raUBP9/swwgjQaXQfFAC1Ov2yQKUCJQNBws
laM9WSjBCClY82qyxpIaRvfmsbbX5Q5gv4RFKVydddtficPLxmcThl7Btgr6OgRbQ0JDib876o6B
paY9pdwuM6KF6C09YYWWU+5hIJuK8i1uqnizN+hx0YvcXlGR19EoPeTw+yschUJK5+ytBIfB7ysB
/AfMvjnkrlZetPmbtkMLH8KVO15s2Uhvvg5LsrgTVfGJQKb/zA7KWEU/fKMB9DY3iBWNpKTj3b5u
L2NS9UDF/P3Qc4g7akiYPjR1VX8qwwbbEYk2yE5qARempOXBpwtTRVtgO5Bs3rune6O3sLlbGfOb
sBnzp2ubxvRqiQDn2hb5t3mtMD3fsbvbNOt0ZTNVOHha6MreU+jwrVtoj++4BF/Kpexb4ue9Q4Jq
nSqwvOw9Fw2wy4Dpu6iZts7en15mTzJtqBdyDl7RpIA6e+JsKd3YemRkgcLzx7yBnZ8Cki0g1Bli
fdT5g0cFGv5XlRaQM2uWn5hKjFE1yKo/Q+DTr/36a4+LmhibNRC4bOUsYCsjJh3oiERDD4rNLdCW
rbvR7UheOX+jtPrjy/f122lpQvQC12hWGWgSp53Dbd6x3y/LrMwzyqALbJrfBcej6PG15GJ3EtU9
kNN7P+a9K1zaoP+LEaDI9lb1Bmbp8zanmYol5KVDjRLQmRfttZ9gjf1j0zRivGjQjmCc/8Fh9wAv
JY6oKyd7y0RsTKjaxT+ViZ+MHRo/YeHKfVuxvoRGrYruc8xR3iu55Z2zyLAYWlFyhYUDqiBMy5lC
bglTGrOtUfMXaQwbMCihLdBkPg7w1yLkSGMgz5iLoLOzuNgkS6ueRPfMWElroCuqnXY2gPPc0UfZ
0YwmBxlaao+swbuThuSyHVVHD3sidDksLNky9ZbSbkpoLvVTSDk8sTZ0EG4MVx54qSltteH0aVdR
T6N0uqk6YYJBkVq7vllpm2MR5zOBRaFwR3ZURnDe/WYySOg7v4OKNgQiQ2SnQE+p26dmdf634Xg7
PO51j7Y30JgFj8Y8Ns9GEgwNvQ75V+E8iqpt6ZwgwWG5OHHJif5QMSn2hYplaZooOaUBp+OGOvbD
1yVzCzhPKpQivkialFEmgXohVPpU9Tn/p4YOa7nyM0uH4e2pIMVXpe+/s4/EwsbDbQfqZVvKIi4z
QbSUnVxdg8ZTDvC4ZxccrJKgL8d3EIG8A+WopIO/dFr4NiRsYuF5jQu2PGFLNcolFEvGeOYy7ACV
gB6i/vjXpVaBiQg3cdEaggeLNY/7ndjhyhdJPe7TJ5VT8SCH+3ueOIswC6dG7CMFL/d/EJQzasY/
MzN5H0nRuJgAUD3eqZsq5K2CHX6LUKTDrdmVgae5A4RwfnH9NF8c2MPtVQQAQKEgHz2LJkTi1opP
uLxAJmmR+GEeCDihWM3QlXZoh2iGzk7kk65rv2oSaB8AbVNe1eyFRVz2G3kH2TavBa6Z9358xljq
GEyNqcYIfGec7gxhEZCNWom4LJ/7TgeMkuDw++EJ/lOmqWdIqtbfBszBxP0M+j6N36BFVP1Ibevi
/Ax/cyUkrixPhSOLZsZcg98ASrX3hawRRTPNhNeQ2Wtx1In1ZDUSGmnl+hBMolFjtPlW9+qKhxET
t+9eVAQvHR/V+AUO0XZ+JT0/S5WPZ0kQCdD5VSch5ghdfbqoUvj7/pTTFiLUz0r0tsCszebZjgfQ
N9YYnKHhGYmhCb4fc+TmlMqIO4cPsLUhBeAfysxqF6gCFgCt4bq0l++8CvEvg8TO3GYH1TjHB76O
0CZlrZdZ4k9S1sncfad37LTaye3g/0vvY1lK7dBtSrmHO0h9R8ADO5BlfXEUhNJ1OhqN5m4CGSK3
EP4Au6hK7c09J0Jc6P1gh9JkzS2OTS/D/4JgWrVJt3Psw/pmN1QsKUMakaXjQpuVEPYR9iwNFGKp
80rkmJ27JobB6mfSlMV8uRg70Qy8IiEnAOmQPZkBZ4ppqDssOM7eUFGNtTKpIAaiwAQhJ2T+vgkE
6q2J4acIfW4sVTofF9GFM87w/zBg07HfpsI6ABtQXvq2TwYdgTzew+d2CMCfZJYjzsKnC9XtayM7
XtHlp1xUUydJfg1kWUmegRWQ1UvhfFbmU3+OD0r1uHQv06aMRWLWQZmxboL3rgHbD+vpmCdLrWHA
sz8ouprgbBLPReVjn99ZEFbBYoAhJZp/yhttXw/8OQ1LEUTq3V7oGQMdYi1kEkxeM16QJIheRdxb
pHKdFdL1WcuGjk2EwgGNL6Af279ovbdoXSxRL/n0Ne6Z4BxArTK+Qk6nmWgupTHnduL7YBJby+YE
aVseZaYk4lk2Yj4uxNCkuabzb+fmO7qVc27NzwYZFqah79CFmjxOItyPLJqqYPMjrIm79KxwpK1l
mIAdGlt6UcsPt3fqdRx7nMZQ94BPjtpFnT/JXndfaR0OKDOld9lfr/9vrOPJqAIfC0qTdnvCoNnP
puVMd1GCXihyT+4PSdUqJ/DBMw0jIF1cy5TIQ6GagZGomWBBDMoHq3QAli2A0hD7LlfkO1jcruyg
mU/SrIGYkvHkDpoBRie7ZMFRk5a/fLdoM7pMTZpVhXyxRIaLT77zArKDQyLUNOqwsJpXl/Cuo2dT
7n21qNP5T/0s12XIe1weiU7xb3KKFzRMn54FGLzla29MQx6fCFQK7GQXW5udhH8CUeVD5h5COpAC
W7uoTbabAVoSeNWpqTZiTsSzhWsO1llBhhIQLfnLmii+pIdWfwW4ooH6ZuAODFmQOHSsZDWo9vZp
obeyWJLCy+B8dzlTVDAQatC279pCBI4iuaNaQw1EpuEv0Zfu1591zRcKs2gRE4N9S+9/9yc/xGiS
lexVe7BP2N+GA5u/PhEMDB0ok/mJUtypnmHaFyJIKjAozTxu4aUwhmHO+pzjKpteIvWMWvzyk2Zu
InxGD1Uty9mr1zLBvQbQ1aR5CFbmiNRnbU3Bx/SkDlRJ9/YM/dFzqq6ZbzWD3HhmNlRR75GiPcai
L4fqwf92K9HNY9icvsLhdSN6YY8hiaT1TLE/qrBNIW+vFn60qCz7xVpeCyqCv/jowUF3a6Lv5aMA
59X5OIQPXKvXw4CzoSdLy5Ss7kMSR48gNTvA1qAtkYPQ0DfmM/G/VHkyVgaOL5NwqoaJKmjEVbd4
DzppvTwYkTtPlUh9HbxnXGKzrXM5ASs3/C+BuMU2QsVQvKc90GAs7Zb0Y9BzSk+BsMwsy9PWkbGy
L7cNEe82v/qnnMkEwkeObo+JfP+5/fujJwJoE5BvcBsVCQbjtZ2g5GEX/c1wSRHlPJWHBz7Osxaw
8V5RtUzBCqhBQcImx+zD7mz3lHJLuQg2hSc8ojC+n6s8Vkau+ax1rlmrcRKYbBTKfEKiFHOqF5Wl
BdMu76BaEzfLDzpM9Qf3N6dMkvPLUUeuUHEiwo48+seVzD/6rUdRffl9uMHuUns420QeDwq5auJc
DZWZ7LJ/ne5gvm+Zrx5aZXEuGeCGaNF0dHK6b77hHxRvtMVTZ1SoW0uKDu7TLUC5DulMHGtrQInX
Rpbdi8mzeCmwTAesWA3f5UF1oS3yIYmPiRuqTxixfBORj3aAqQnFL38xJtoFOXvb3M7Pg9BHo4+1
5071nVHL7qTv74wQeHbZ6DwDfxhmY45FIwIpuXGP3smI3wtvS4HOrIq0wT1e5NkEwkWcqQiUUCE+
FtaePRh+nD1oAAeST0dH3iVsd4tNxyXFTxgXhZrUSJRF0/zeCgGrEI088TrrSpa9euDnz6TxYK/s
wesaW72ZBvLJcoBos5u6hRdxNNAh6qC3dNPFnmFvy/SfffeNm0FUnrpDm0FXQ52k0MTit+aH3a5u
1s+XOZh6qhmt1m7pW1FVpLSPJ/QpreNlYwqeBUGUloPW9LQZdOWWjE13WDpVIbIjqJXcY2iqDMAF
bZkDj6pAqWdrL/POUjTZBGvYErMDZiPkUDJtor7bNqkXOBez+UOe4AHY1lM7i2vZYGiBOOdHUNt+
RkEV/2EEnnu/r6FI8Jw+6KglDe4jHJqWuZDxDpk4HDMW07pcT0+FHCfarQg8xV6fNL+4QrNZFlex
QQawiS/SMzhRvxmw6+ifB4JGTTdhcQ3cpic25FaMZgmz0y1t45wb+xdubctrQVRQZQn0SuEt5Fj8
HGy7leWaldawfnrXVtpzyA9yFqeArGIlaq26aJL0DW4Zq4jGU3eNdso8VDTBcUl1r6B7q4eM/zUr
XaJGgza7zlTLe2IhpogDuqomuZYDvkHrsRjG1DrVU71iAHueLhYw5QWajbSuvQ476+y2soGUnT54
gctAvABD1xWXt6xmxuwnkThbOArxhSgoNzaqSjfxld6EIuylmZf7w8Fc8hbeCueCS0W/+rDJE3il
ZnSyHjRdtk9wr9mObBZF9c+4WLxzUH5AJS6bczUn9BoqqYE5xmDez4Zv3RaBIUGg9geq2tSbF9y7
maeXWVFdmta/ptTV3RNVYBC+m6+uLQlH7JNOJlY1n95x1VnKbiF5u4W8cAukPi5kUxXaDMsVoXww
LhaVe26VR6oRuDpx96qEeTi99lUUkEIL4CbMDdMfHgxB9WLylzwgBn+1ElSm8dWpedjbgNujgYXr
Mkyv1yLRZEFiY4gP9Zm6bV2PZQuvBRm92fLtakcyvNC9+t5MsHeHhXCCvIH/vgIDeaDN/IZp239q
u8Wrtg7XaGfs+QBPAxy/6TlSG9AFQWyEQesi0ig9zd+dqXqrv63+sZ2TyEuuQh5O21ckA7CkJ2Pa
Lo+2sFJgSdR9rY6Ky3gvTl8TjzkxX8t7wYcK0ZMQ1MZWDs4OaQdovopoN/QhetDtRzK+sAhQPc64
XZXa66j2N7jomL6e23XMCcwITXTuo7kAXsjRSBeEpFWWEBIgiGcQOY3wQJnSAJFrw98qC94mm/59
KBUCoOuoXx0GJ8zUijr5B+987ia5diBoFROl4EiFi3dG36T3ghoSN6vnTNTQDHyYkHwxx/XvEcyf
n2E04yySMxL9wVusrwAm5E18yFBIXb0H/g4v7uetoTJW+z95DStwImZKbxx9xOjp9IEZcHCiDm5X
dF0FiQqcnIt9JUITOz7GykRhDOFPWEaEEmNmSwN3v/lR853Cl6XstZY0pcPgULnaWNfD+Cfw8QGP
hJqUfAsil4/u6GP62INKUQZ8sE2ClnWYF60KwHG8IdzzFMhGcWewIfQlvMqIbgqQ94h/8R4+q57j
4TPM/mBATuZYj9cUJeCnhLeCouz+IJBinHPvooR+dRTBthEHRHN1ysi2lxbumS0s1YgMCxmQ2XIJ
prq2iaOYrnzYIyC61MnEdz7x7lNA80D5vhDvzaQYu/omjuF//qumb7ao3gbMcJTzS/6ACI9BpEKC
+83ZLV18qHkjIBYoxlW4+WNf0fuWAvYfuxQSqfYYnr9EH8TvQF1fiJxmDcWU6BlDJBaPm6TGOD3i
cpxo7YsSosc6LBSe2oPTUIJK0fJ4RzlUixxwLav3YvnKpFDIr0bI8kV2CPoKWULlYrL89SaQOmdz
SKEMiqLK8Wf47ckkeOGzhEJKcg6cA8fcfkVmeKw6pRxnhNPOqarR+3ThjpaKlE0b+AT9h70RtC11
4Ap3ip+hXZ6SYHJlp3f8sHpBCivMwPVaw7no9FtJ2FkOM6M2+MYXHU8IKa2Oz3tnAYsEzCpYV0sX
lF+e+Z6KhasBATslDsJtL+8y6qWHCAnjmq5cTU1AXlkWU2K/GSDpkkB39de91Cyq3OpCMH+UPoET
JCIApTI3AE3KoI+//a800BEGbZ8YMifv/JSsoSFX8HiiY7sKH37gwxI9i3c6B9ltPeFpzrw51Jkd
EZZSwF2cUrtRfzRvtbJsJoXuSbokSNrzNmfS2W/iwy9j2cCWeHOP8el0Jvw7iUMVnr/UWeCWDRc7
hx13nhrSdp4FM3L8jnjKesdUowLm+X3vxkWQ0dtFEFn5voqDvx8TDmfaqHgfKRoZdX0dL2Y12HSa
xoFvJo28mHE/DqhgbYAutiZT79u8kSyfz9F9e15c8+YGzLXOMGuGjno8GCdufUPQ/a63Sf13OIfq
h3iILhwN+LcOTOTNTi+odgOrMI0mN6NiHI73EJr40ErsXVQ+TPforUIcnLl/i6WtYhr6qQDj0IY9
IemZ6TwUfJpRmqrbtHCigg+UjDiNjKwie0EIBFk7j5U4ylPuLOEy7ubKYVieLJw2mkZo4GJZjDN7
NHNL8ucTk1QnnMZLvv9jyxlodjUAQnrLT2r3vIZIzH8vUDMBhspDqbiOZIZnHFFU3UcPJGeHCW/u
NpzdlPVBI1Vh4EDz+wrP9F5LAS0nONKNGSvXl95/V2wyYl0URFNP6lK1hrwV+C0mg45w8Jwx/wIK
5PvhH4Uwc1pV/bgwSZyCZI2V9hvMLl7IABtYKp+xaTCszqwRSpbpoLIfBV7kNfhQocUYt6WsXajL
CI8BHd91nHLqMVC245HgebDf9f8bbIqMd9KucQJAo01Sd10X/WxSvigbAFPV65qcRXC+H8f5d0PY
Do2gUAY6GgD5FXpzQtKg5JymGJr9KFZh/jbz7eHGtyoO5EkW++CGyuCJGPp4YpGCqr3ybhVnTz/7
btsGbRivGNOr254I8/CW/uyUbMGYJSyVx2SAKIIgrZSZ02LXkaVlGVSMeIW66IW/V9RHGep9AH2q
Yj89Sj4zAxjjTP4a6fY4SG9+YWjYss3dEIKpRHf/llE6rzaETDq3UYGbEBhyoCA5I1PEQ3cxZiVS
zXdmsKxKVPrrnnbs1jrTyr+OrLwF1s7Aa2o22QFa8gzmRxJtqzvLwK6HaWzNt2C/cpdmCXTDVJsZ
RZoY0DcEpMELbOeEicpzbX5GSm0EAtIC6cZe1pzgeP3UozvHQx0Obwn0eHk0Y1ZTWdh7QIWKJose
DjI5Yw56hEUF3I7uqzwUufjkcZPI5Nwnp5x1t+abj77MmZrrXkZCj2xDJmN0iUs+PEPXdTSIfY8x
vdy3x+yG2PXV+x3SOzJ9VSOdt7PMW4W2ztRo84BYZf8DfkvN6ifa8yNEl5QrgWWAScinLhJjKqSE
TSf9tR0XsvZyRSOm6uCMzXh4WhzZaT1McLd52TEIsFbJE7lsB/Pcp9bSZ5rINg7Xb/foAzQ90rUo
YRuI+k1naRGvNdW1IfZTCih2LWqod1SzCvvCAbftTHNxHsbct9d3+IPExn1909ID/tM7Lx5J6krY
VrFmsyvajOd7L+UV7h1RwZZ6hm2qy/BY/HzFMVG9SogMWTYOHFFXzIy28/iMyhUcK4KemtK+5IRJ
QmxZchDnGZuwroWq/QepAfMvdVD2gXguxkStkEzzlo9+uGYEVQoTtOKw5M/YcMRM5Rx2EFMz/MbB
CthGWnB8OOdINDsvNQuOz/kC0CxvpAkVpoKOGGCgThqL35fffkZstTkrPfwz3AN2bIJqZnawGJDF
QwUxQmp/Rf/S3odPsReAG/LQ4xfogFE0MVz5prBsT5lnarqqo0iWlsnCaUqZ3GK/sc8tjSH11+D/
+2qGE44xaSZMzUVBwOTdg8VkmBxpTUjMB+U24/hxiSHHwD5Vxeq5yCaAsAXyHGdVAfHSdnzlqFZF
a/aCDRnBc5Z0YkcA3Mhyn92OTuHiCTvK88b8fI97lp23Yg+aSZcQmOo+wKzaTHx6ccAC5cmU8C89
jKRY5/LNcAAj0N/cr5PmvR4DYbc/YpZ6FquIKvN6S/nW0z+1pNKjYrCLEjzuDKgkTlCBwZBuWYoX
L6zYI4/wik3fzyb/mDunzexzwQNutH2OOA32rvzOa4D7jWiA2Im3CjtpzMF8xlOan0lnMHPVZJ6d
V7GZg6sm235sE845NJOrZ+lKryQ+qoCLO4KlZsmm38tOk0ENeIAiDl0IdNAI/yZAAofpET9SnnCi
8St3JfNFpiXREMNlS2rB/mNQJGgMs9e6rHvrszxfWTcd4UiWEAe/Uo6rvqQRF8BcUG+LPnilB0vt
ymi9IicB0H10Ur79DlU22uMlQJXxfxlh/MAvyjrO8oTqW2H5e4XynnjpBv3YyogYdu3FFtUqgWzf
chzPEGDpe4I9AX4aOU4pJ5ffLDCWT2n+/LNtI8oyKjO4C+/PKbLm4sSCxDStIjpS1iZILHiuecdY
TtvPw0ZgtXrm1RWZKc/HQ9Ay66W73FaV+oB9JH64ItqiBz1xx4srnYiaf+K4WqR46K7Uec0MZtJQ
CmP5w/UCnypmhZuONbbCVnI8q/KPk/3QGiq3zOaRf6WvjjLJM4MpEvoPmyOZ1WfMdE0ZatdQl0Q6
4YxDt/EUqHBix8+Vt9etUSnvAIJWvhZayASXzBR8FQ6+Kz4LOhQd9VPTMmolN8j5l5xd4Wdot3/v
TBlmt6FJyHRjtQeK4rgfaLvjGKACRkfYcw2jZZQ98FH5zTQtIvd/XslKoWrixGnA52wV1jsCH70R
ibjJxP4gYGodIkk7aIwqCOejDIoKXO7t9UDJlDrDbmHpHSYiCRFskJ7e6XXD4IO+JcgGVI34t+dR
mo0J6FJ62XCan9C8Yt1TEPkAJxPgqnTkRoE7/84HA9ABtLJh3f4VoAMzvkYHdm0cuJ9br4ayLxJx
oKmrLMpdCOEmEg9uV92A8fzE7H4n2eSyfCxaNjndtZ+IC6HlLSuQYRsdSzcU9G6om0Xp7BNJV5wj
AJOyCfs+fktTeiIc0GQhlP6vMQOufFuvCPb4jj5cOMaK5YFPDjXkj4xqPYJFfxdSqdXeucsmpoGI
Z7wMfKkYWlM/1SxjS1CjmCOlAnS0rS37AOpq2J9I9XlfUMaC1O2SxWzKHnPTQr2b2KA7JISgcg5p
VuF4rLaSR+/2BrJHW0kWFvzgwUFpwX6JAqS/6L3ZFwGNrvfhoO+KbaVGfiU20+TjVRbJsC1jWMjb
GEt7meyrv01YAckALMkakZrw3rS629hpM7Fxp6pxjDu4glkozhAxllHKbBWVmOHts9pJT7hz6Lz0
iMtctL6KTt0GFJIoeJyePLiiomMpVQpu/Nw1dE4WwwUouDWlXH07lL85peeA0+9QmvhZDCHBy+TW
LIQvb5of3RQGt3af/DGCt9Hr0G8FErqVN0SrepoYucd9ibKfVLspKE2BuSA2v2Q+L+ZtNspBI1sE
1+uARxwsdXSbPWNa2rUIDqgC6GTOQwATxbYyOMFd3p/cRJnOV6ZmOYFiq1AZc3RuNCRf3oK4rTqy
xcZtqf2SzSksaS+0G6G2EaauKpelIrYyz9WbN1+jRzBIimKk/9g+qCKz6vtRm+eUr55IhoymJ86q
rsxt5HT8B6q1mSQ1NVMpDCQNw+AhofG0NEmeAdmyjTTs7eOjLc4rL7azyFvS5rU03uKr6a5QjG6t
0dJxf1ZiHYj6fW9VpaI5FfDEBzKCmOYxpso1v72P7mYohRqEtA9fxcAaM8RU6mdQzqnPTm+oZE7S
QKTd21p2NnXPkAADpPaBuWIOmFQzfveyIAw8JobVS3jm7fE8YMzG3PRnJllLve3a/1Smsg2+s3Cc
r0IU9Rfy7jVJas95fLMcCzSCyBe3pHQFbyrA2nJkHi5CzvXO2Ad2r2oOTHqamv2NZTMBoxL8qslR
fyvu0o5/tTjJ+gOp95gF3xJVzg3Tj1fFpPR0HIyclRN98KjSiVe7JTIYYLE8+mD+g4lxsw0Sdy3j
dqPVPYzEHU4oXZJDazOocGMIGfkUw+gCgpuuXvQv1ANR/ietkhkNjC+Zws13K43kCUCPg0UVGTHh
FVYylKWvuj/2iWLI79P5HIcbZzU3sPRfstWIYFLUJEstUvOad2m31d28O3ohGNiNByCHeFfb8/MN
54wVFug65eg9B6elMrjnPCQrfzSEt+O66/gYxpc/Lngg3JqPCnIZ+CyTgRk4S2uvnNjaBEbPfeTI
xpYaolCdmTZpt3uK+G2MBTq7pJFQ5RdpSYm7yK3Xh7W/lvOTI+pWsK4wECxoYd1/gbFXY10Au0Y+
5j76OFyzaCOGLgaXmcE53+vOKxDZZm/viI2+GrskFkxMghXt53g4A5RmHR0BFZJWCHAxlzj+gTft
hsFLfs355OBNeh2lpEcqNPOCdqbaZjwYlPQ/hX2PiLVFE5elp8NPiVYKEqAL7dr0AePKDWmjnI9Y
3bLgssmcE8eqHdO3Cx5ApePYmQO2VEE+9Mi/A3QJS6EbrqcgnRSP3lbXqBRQj07B0tqryRzNr0vS
SsNqGnwrolDCF5I4PJJqNayNipdV8uwWN6dvq3JGGb8jBotXTsamFJFuzX51FZZ7e0Zy3FcFSxBw
9A3VvTCGi7l5oMefjBi+Oynoua0JYghICcBAGIy2cirVL7SMOpg24SujUvSClfYcLJfAZ7euw9Rh
91sA80JB2nDhbj1UFK4x8clhtTTnCKfi1dZyYlQi9SXyeCGAOEVJaJLpWcb+NNktFjFvT0AvfU/p
CiNKTaagNcgjBJI9YIFJHcZadJgOs3/um+doWIDD13BZNehxjNcpuc8ZK2iWz08YoTALstn/9kcP
yGpjTkfjhYcxb82or9iwm8cuxn3I80VlObU18C3gWE4Bjl75yhIHnrsK7ZyQb13go+KZ6Fiu3zhK
gpLlOGNBZO/lXo69R4D/sv9nvasRW+Bh2XlCI15ZBiAZYOyZsJD9NntJE8ctT7Ah7S+Cgy+EcbS/
vjoAOtMwCWrzF7Tzzi5KmNCE7Lv0WqqEWmOvHml/pipvv3F/GzDtp5pnnyDRhsoXNrkYW6RFz/5Y
m3+j3y8sHUUdgk1g69LkijjnJEA1NJ3VD/rzMA4sKvEBeCvWUMQ2Jgcu6SiPQsOrrF9Lkkb1i0xC
2bbT0GJRSEsRPGgu5t8x9zyPlM0M1neZhrOx0RHUfEIGo++n8IG6iJHHZR0nBLsglhC2sex9OWED
NDQ4JuVKTqEiXD81+7DdlYnTlNu9pBPr8gfuzqCq/SLZwu2dDCuewVaUzRghW3wcTWKNR4lsm56H
izvn3n2x+ovX/dP/Ru9Dq92w2SJC6rWgnnFNCcdCqL7iI7RZ/UgvNC2S1HL0YEAfjTWQVRhYQxUm
vK7boV8odT9SpGKaIcUt3AdhiVCVpd/jdq+y1PLC6173Z30DBT7Jhew6OXxQ33UAf0JE0PGQ7bei
zgQn5OxnXIZCtgxyc1paUumY3IaN/N/facImKC/Wls4bugcVXJo5CV/DzFz/x7hucBwWcTKvXpjb
3NMDdeYQRzltv4USAu338uP+CzkFv6jxfJUTIAFDqV4Ivg9LVDDwBvd2FUczokaGUjg9taN31VlA
nDkHs1C12kVdeg7/GutiaJOf3TWZt0jZBAC0sg97QcIyoX0Tdds01CPuYkrvCS5Z3Ie6WLniXcet
WAlrAmJUQP+Ajh0v9SHfLKrlQ5NkltNM+HCMrVIn+5VFJoxBqP0oRRW4btJcQpEt15L3/2pk/cxE
Cq5tumbtCL8u1GwMc1Bb8+eBaprT5D8lBrwVKfeNFFFe+tzD3iSsS4ZrBuUAnPEEIqKyba5wejC4
0DpIb7kHg2npzkrvfkO9oehmeeQCTEhqIC2tm8IaBoEtFRruB8f4bMRUg4uCERZaPH5xO5bqbGv4
0t2EzTr3ej/HIcHVxGMbw+Y7CAxQw7FqLMRkYECbeWygUOCGeaU1dsC4FGOiKHJiLJco9m2Vlnvc
WUpaZi7sg6T36mUjPcar/24q2aQ8VRFbQb5SOJCUsO3lpj+rlMeEPjGR4uF9WTWlgZq6R8C375rr
JVfTd++iecvP4I1bTmTr/GH5POTrEJSErEm+UnOSOIhW62yB6gyMvUGVrJngTJaca0qo9y/E2FwH
hhQAoXNu2kHX7x70lt3iUj6StZXuEbdIEZQgZBlJ5HlRrVhbYYhPkNR+sOhEKb6ffIeIieQ7caPx
HikgBtTfGo7zFprvPq3a7tCnYRQNhK0ug1TYxq4ZnFisqepfI4Hdn8ZHNGbIOZff+x/h8w5gCZFr
SfUVh2ksbsbWqja85Ob/9sCpews6xlQHo6NNhzzxYE2q6myaPpTV/DVsx1vVsxeb6W8ht8ql5sxS
kwY6mkReN4CSQKGXoiK++DgDGqdyc+IMMDkeM1lexPBY3RPhhdCLaPdcDNxxt6jPsBfJr2Pte4J7
1jWI+PPGdAGY09QbYoo2v03ueBeGkgUkrs/jfXU9uen4D/Q1ETPhRmw2gd4v/8yVU08BuxcuVEcW
MBoOU+ugV/ezQ7Ljf8SDU+PQVkFkmMy6HQPZnJ5DVgKrhwXpzwUXTAfrKQshAMjP4JovF8CKca50
I6A0TRnGlfQI1SSUjNj0jxa+5TFtuMD9glCBqPTZdBzBbYLVYA69JlCTRZpcB8Y2Ygn3iOlYDAzk
cSZpRv/yv+Xn78iaDRM4Slv8/pLlPTtX0877k9pOJjqXnpiotXKHe3iqIXv2od2GEKhXQS7k9T3P
AnF63t05qyeC5grU3QTwpqzHz6LgXCkx8q22bOPmhx+3qLKES18ZVGm7Zn5fal5Vs/95TBMQ7Eq0
+1EsU95A5T6MoNX8PUSVZVuy7HzAM9xHmmzmGDcMRNmQvEIlXCSP8pc/TQxUyc8DCu4eVZEukSnn
Tkztr/YWjNOn+8/8+j/RG4aQ10rLRqlIPR/RACRh0xbUetFFzp7yHvEchGvpI9KZNOF7a02XUsU+
yfH9yvN+BVpfb5DUZltroyBmBzajv2i4vmQqy0wF+ioyb2D8uFdK6RbRrfPpoO3A31DYQgCDgLRW
DQgTLgTZGLWzkM3hIpwcllfR/Ll1BFcwZAYye4c70nBItxxPhsxE3lS4rKW/vC9Th7ZZIGVIpLXb
YNknV3hM8RgwS6eNust0b3hX4RMUx1royV6Od21WY7QjXUlcd/nYtUU0tMg80n4egK0FCUdHeKEj
YNFOVJWiHgyCeq8p1olMJ838NKv6G1rp+KuwE2+KUJ/ZLJq5dWmQEWn5v3ArWcNVlQjLp7RpJgG5
f+c/1uISn978gzfC0/axOPrpGDKZZdXsiyM6oMeSMlGsn6iTSj7fY4Gmlty/5uyubHMfYi9fmwnv
fDMw590WQm8w2qCvYFWmFVo0FxGaNndxi1ZFrmH8M83O3TYmjpxqKlD0aqY/fX4Q4bc5Y9/W4/jT
5Me3bpsR7njUVUy1x1TNCzq90Yq5v8gbk0/hY7A3pDl5Q0TEE+0x7L8t8wwTPCr0sV7dFh6yALDT
n710WyzZsiSNvSqXizkwGwmdUwpXDSckTru9aDKdHIhYSF85tkgXtQPn2WqqFHDqyUWUm4e89A+w
2scw5lPbGLVHexg6ULA1LoGPdCvfB3BEUKL2tLEu4e7F5lHCPPZeTs/NTc3LGXyIiwfbdcibTBiV
NB+AVth0MN7pWXbkcpMPnaeqq4CGZqRwPEYzCo5d6FXksXPjG/xZMYeVH4KOx/kR7z69kZl33nGr
TEHNdDnIpQCM3JQe/JrITAT0J/hbst8oHSTgBZtiMN8+KVALh1lA767atfoOuZajFeQ/J9uyjtig
e78Ey/bhMzDCbJ6BfCyh7QipOXucdvJ2nrJSNRDG64aoKJlPpx1YQpOf//6blQ3MQ7C09fVeW9Vs
oPqzaa5Nr02xrNkyVMKfbrQV+ridKnNNOZGGOzXTjQBSOYfazsb6c1HpMAiEYh17lsGhiVf3/ecU
uELo0ARc4NM5QWyF+3DWy3216U/6JSoQsMsArc5A+B/221sxfWGnAPvELr7/B3KIYiTFY4QZ0zzO
xSAbdcAsDg8lNtYbGEq9RtIDQtgl6p8WSdFrz9bukZfkBNQmwz72VoJZBS7rdEzfwYXbSLtNRIPm
9ai0QrZbyqedUe2uVwMcSvKMunOTEvWxPMKnNUz/gZ+8Nuszt0w6QXJbzYO04SJ55s8TefCY1NYa
sSZjEJRe1XUymakSuHF/jqDvBa/lHuRJmwHdTGvoElyopOIrohbC5UQydSLQEqmW8AoQ54Jrg9aV
UjIpK8oWLk/7UBnTO2KGl3sedWKcm162YRGvj8biUCb/vJrw/NKT8FrWTKZGkGtsL1hk8hXTN/oV
NDkIwy7UPtK6NpwWGmJmpUm4Ysvi7Got87h9c3O1OQiwLrdHETvtKqdPumNqy2l4Plr3U4/qTkp9
0ZkBNpOwXKUXSUeaJfjK2v2KAPJqdn9KkyLSGTNSw0t5eptbMqKDp7w/JAtlRCnKoJr49VtxXNOR
zD5k/gvMTYqNVae0QprLGQxF929Pvg7eUS4/qKkdQ6XMLjjMGZE2iZrKdr9iML6g56ST/nVdEHN0
cdAg3QW8L4OWSqQQvVaSfPLI6PfCsCr1lvoWR6sPZ5f3HxArGA2GOnB7M7zXVhhSoiboKD2+km06
0+5vafZWf6gxUHZoRvJ+SAfPIbHlX8FhTrcsepeuB0rzFllBdWJ3WO1K/KbCpPE/K4MmHecZEd5y
G4z7CpAaQri94bOkHl3TwZU3wXvBKrB+4Qv6QRcZmVoUvebnqmYkRSBs5x3l0G/XMWYpL6SYZ37W
P3h7sm9NOJmOXaj8R/S9F2T+yFTLrn/JoAPBvUWLr6AaA3VS25ix15Q5gPkXmmvOOPxz1rF9VRVb
bmEDnuknmUUbH7yPaFgfacwW3AcRxkPGVrz4fEqnSJUzwFPdOWAJXxVYghfqZsXSA44iAzRSXHuJ
2VTXlDITsowcDKvYb8f+0PytfqJwjtCG/c2LFqCw4yhcoHmP4T5ikLD4vwCoE4iL//AdVuUYBQZC
35BsQc+OO8RqE9Gj9FvRBcaDt/kSpF8HM2HZBueSwnyYJhrlh2kwo8JJsISe1SmMzTbhykZUPLU6
FICSjjCgDvKMAUzZdOkbGZWfmbjoRjoUOd4cig8M0+6OGq5fOgf5hAcDR6Panw8FzqbGayDggQTo
dofX9GC+ete+j6oaHTqiJtfnGSZ5+HsjVWo4lrmtpBO5dXoaSSk18Hl+KhDy8LXqYW+4rJR3Axo4
5yhNVYEQm5Pm1t0Pf+DX4aS81ZAf/KhXnRnR8gjhRf2ncRktlz89as1teFJlnRl2rAJL7fc5SoSe
plvJuSFvyyBlU8ZodsYPSI/7OnVd0Doz37gV24aznY5lJ7HOuJrs/m06IeahCWgr/3boV7fjpqWn
zKy3oLj6VdrTwcIkElxztQjtEE/i8R0ATFXBzTgDjzgjtSts8osQWwU2zfHeUD7FDz5tabyE3pRe
rdvcpHIDJS+L7PfPGAjoVQyPKWSskTOt8ruaEkHKQnMxqkA3rLDcNIoXyJxlzu4NCzsdITUiL9nP
Ao/NqhNIbLd/BCZc+yF9Px4TMZcO+bWYDBuMuNmhfv/j0Vad1UqlMO/rYIsR8Tua9o8OIGHXhC29
leqFK4YdeOysOixR+KZ6/xDW1yh18AxgUgroYjfbgo98bL9aXx720Vc2/HWDscdZjDso03Rm8Vyg
eEoVGqYehDtVFpopocs96RttLz9W7r/S1s83xQxbSgc6xVQdbxkqfJ84NUS9sRIb+3lZ/l7HfGzE
nUEps2aNu7idbbzV/ls6MmeYfStLd7EfZEayTo9zXamQYKztKTD6l+DZWcZEX7Zi1VsTBtAk6fj/
V/2aau264k5MD/FCrecpv1jDaZsZyoILnAnrR+n20PBJlxcolMvyYCEfD1VA5oj2I35MKhtrIk7B
1lRcVsjiSUvBEXqDHyo7RtKDLpdyKT4nhemC2NVFBkPEI2J2fqCHyxiSemsrQP6zoo9Y7Tpl554r
6PFxACwV5yDVyJml/A9xJcUGrmkAMud6mNMbWY5DGxp3PLZaR8ysGljUpX8zeZqVly+8z/qAfuFD
/xZVZxP4G1WdO/ys49Ossf8YlVbCMrh5D13aKzRwHYt4JaEP9b+npxsL3ygRGwrfgcLWm56smkyE
60Nweqpot9somP0BIU9bLA99rIPif5rvsNhqa4tEominlPkBFiLT8h0ycrpbDTBIrOijQk23N0NH
FCR12pFHEMjwC15BxHVDess7avslGPncugjS9VQXw8gczB8/poeejZewHHD8zqYr0Uwy9UbIGzDP
Xczwep4PVWPi3soMFI7hUZzZW82qOlxoQhMc/e1uhgIZsXiUW/1z3xU9DhGTeufydGFveG4f8/+O
bu+k5yxnyLzvXEDIHy1aKHmTdq/JSQjnHtqoVGxBAGm7SLe6tEeabE+RVgngIzTObY77D6VN7J9F
/sS1XSxaHxbe2O/4rkZgG5iXbNOeWR7FjWQF6z2arniHLvBL19YianSH4j3ZEFOdn9aRevquAmdn
j9YuUnNGJf4rnzmp8kg98DuZdK9CLp2PVQbcfs1O4+ETvOl8iZcMaFOsO0EhZ/MG1/r6wiXucce2
ggSj91Z+hBpMEFtTil1Rcrcj/v5vRc49xGMup+wFZ7uC8bGwiCwizFDXzGh22C8qD/PtIpZcuYj7
m4dhfV8hPTqPW1fND11TpTdMgHs2YzLzsDjrlVg6A/aExqpAK8fI2VcMdHdO9E2HCl4tKoXMQzN7
zHR64WxLbj4inqhC0S4aaWHlJPwcTkxT5pnUV9UeZ/GaZqfAg5RloLX5/SD5MZEW0UTb5fHUP10k
GAvl6Z53qrbpzQ53t3Wbh9aMQn8Z+SqM0+oslC4OYKA3OEG7oGLxuGZkEcyvGU8792xIsX2voRQ4
sU5nJRkaudWlbGT/QEXkHtoXk9LvYZ/k9MNCE5ViGPn3mQBqkXZLY6bbZfH+uPxnZYcaXLVFKuCv
PaRmdmhzI+ukYfh8Lamo0g+auOpTAxzL1uwFm9POfDagfVcsoQhdM1s3PrTd6Up05T9ndzBNbTMO
ybQOLmZyVU98d1PR+wMxmefP1mZhika0WVJsZ9qzMGhCNd+rcno0EOzDvKuG7qk3jfTTesmOhs7V
58WYI4K7MxrTbn48bwAUmxkKGk/bw1EUcwHN2PdB9nst6yvHAweCcNZ33FXmKd1y/LoJwzG3wKma
jBhOX/o9Q483Qv4ORcd9eeqfjScNFLPKJbAH1HSZBOoEGYeBi/J7twuoN5DAc3XM7rypp33cdVKa
dxXZetK9rcNejU1rrZhT6o1jrge0Tw9QwVqI8gWQYW5Flab5WctXDwY3LPwtqsOWUCDTY5dXeSfv
QxCSjNDvRx3HB4xDwUFsScClQZoY/Yb7UM2hkNWgOka1JlgG4AcImqKBIOZ40VLI+bFRxqHbBc2q
CApVC798oPk+74EB8tZ1Ak43nA2G50p5fzobBcT8Ia2YYj0ST663IkDEGIJ+ysuwUGxQsuPVdHKW
DJqzj8wHYDDCQgY3e6HWZpRnxPdPcG3SU/DuyOxkSWM4roY0bgIsw60TVXhNxfHwt9KEyPcl+3Lz
+Q001UUjxUY7Nk99SheFZJAGg3GTV9j92karpaKk+sJ+0cvi1sjBhgwM3qsMMKJ42S2nzfhLmumj
8qHZ2l3jRutwzi3g08C6rZ+VRNQA15tDj78ESFnVYc17bHJIKMJifz2es2vE0aGPhdPv8DPlm/yq
upml+Kkos5p+NIs0RwSmlcOoy4XVwUlYv05s3T8J2ew8mKNyP75JICb1z6fODK2pDN1PlICZiWWw
TS6tfgkH5pUCanLam0wmBeOq2GlxMkyn+8YKFsDgAH1M0/pXOy9u8kZJ7nN7YOgI4SJV96b9aQb/
pVRxMFF//l2vze+uM3v7KSJQgII1xnnNj8C4F4kYorPPGsjfJ/uWnVKnVkeOTBsbnScyZBScKS/Q
xEfy2KcnLpX4TeiSILe7sfP38VNkEfnvvqeUIiuHBmWdjE/6rohV8UE1rIpovXm0sFoHgf/XW/0m
1ynlzChdk1dh5mP/3JrnVDxjVH0veckxmhrVM20zhVL2H2F/m0zu/ssJ0QoNme3p+EP/3s8GsHTg
sQo6A77fjXrSHAIYpVVR/EJXTcEXQfsx2aZnxc3EK0RscFk4nMXyr4kPL0QqZYH4cVWwFY3YS6oi
jYI3TCy7QV+pLI0AWAIyzn83/Bjn40O0JM/xBRktqoD8yJdWoCWKtifMeZ3UHwMNIWpSTQ4muI61
0kO8NCk1o0JhgvPQTh2H68Z7iMh+12Xs2pRac/csv8G9++n77LDgh1LX9K2kWqoyplzc0Q+06r5l
bhuCs45DZAhv4AcIAJrPdGNKpzlb1MXf92JsXclw1p2M0EJ1s+pNi4PCo3c5NaXfgnb1l/81j0I/
g5qVPfRW4ZBUBwwF/k9x5N4g6YDjMg0hptlHpTaPFh67WVKkN6f8BCcF5uvI0Kmjrb+ptLuCAutF
Z7f3MjomXH1BCDI09hWUdfMp9Izz1u8vrva8oZiK7A5oyT7SNht+Dh1B0mptKLG3vrubeWRcldN6
9PY5S6S/xnXNgNs4KS+HSq1OuLLEmkzZxvtSSPc90bhZPgLOMKBLMu76tmZdIEgAvpp/u2N54R2/
VeJNoB5uFCdfpnC2O+oizmV2vRRTF+SjK2Uh7ZeBj1mesJosDoEq8eNcbvFA9LdcFggOTgNhh5cT
CavUrrL1fF0xSIpEWhzSbp938/ttPcR+h3xuAf6v8olDH+MemJOn14xkXTpSxDzS5LXSz7LTl/do
e/s+eUmHtCzxrUE6bqSsdvBDv00be8XOf09tB/9xpAA/icjTVS3pTUgfDKBhaSAjpPm53lkjdOrw
EyIhaOyWymbHWMGiGnJS3B9zkCUUMFFnFu3ug3Rs4Je2CDm+mnzbPOjl+z6E6muxzgm1NDM+CMzq
NRhe9CsTjzPYsRBO8mknVtH3ar29oxViaHvN92earVdqoYY/wFauIfpKkPxJJ+ar1BkLj0MFWExw
GJ07IVX+Rbz1szHE2ZkJVfRDip9rNA+GJVXzBN1kVMDM8c+6FhgCj1hMhsCt3Zd5iC2DQs6ascst
P5Qwl60/TgahkxL7A43oW2QG0ahvhk8DNHxxIDiv35N1sFdWMklfWwkbKNidJoBmHz+b65py7lxP
WDVI1dGPLkamdXFWPyh8quBLP+N0/tIMV22UkLlNAno/BVfC11eIiChUm8ZaDQ3NemvK0YEkJLLk
/ZiEq8AW3jyGHc08PFar5uRiFvIp/kgBinpbsfuDCieSer969NrHgf3cm5YGU+7sy/zn0tYHoCYP
ZtnMqMy5nVdyXNVp5a0LjBQAi6GIS7k+Aan/EFF7ijgRyCVA3q5y/5+q64LrqasCCp+w0MxMJ5Fj
KvvEJ+9mC0zLRCtTClNNsVtmyzXw2iw8gOu51TAFHwOP1CKUcTioE/sH6Pb61Yv9KOoGxA9S5w8I
ONtC9Roz0aY+Qi16hKx43/T2asLWOk9h/K9rCaCI7+xg0293Zseb5wlJyi/TlIVO5tE9tfSiX3CE
RjpA50WuS7H5CUoTRUpVf8AGVumt7+2EkPAyFKHhQCxkSyrNcIM/9g66Yj2oXTVf3edwVVoix0hB
vQkatetBb2llXd0aILClO3VXSn0CY9K0o7hiDdIM0Sj7OfKEzjINmK2vrVVGmRuMaR4DBqDSJSDB
w1aYFKVQu0WGU3PTqu0IuGVX4fpBvKSdKzs3jVJGfPjVbkGZGnWSbir0v7wCwnaxDIyE7LHHRfFN
jzDsL9zWcyUiMcuA6KQ+ZmoZOqqSaf7LZ7I7tP35KRPaKB120jgmKWSnpM7eccB1ONvSQ4x2B9CT
475zNEk+n6z20YLwqsHm5mI83/Fi39kQrddP0IMx9fSG6H0FU41v3J66Jc9x+ZDUjIMxn7eOeak8
OWSUvD3Msw8gm61qA0wMRr6kPw7TQ7wWHolzxuNkFbLoUaGq+8rRsEYsDF+gMoteP1d2uknCXJZ+
NuW3JvFJOKB0NxiVWGv80jQa63SSxymNQ2DAVAtu+soGAMdwc2C2ZbNAIU5ysRirAal/Ft3Uavcv
YalThhyisjc4YA1muPdyvA6zgrU9HJI6HHL6Cl1WTAOK8VAwhBdiiJGIbTJxg7BweaqXlh7A7Npc
4j8V8OPQkGY2wCNy85/MmS+dkPc/zNR20N2sTo8INXFyMj8/sU3CtFe66TQwXm7z+DZtd3RdhYcX
d3XDwHEZdwpJJ6e9dTe/R1JatKzScSUYzcXh/mo9FPEVLB9qkOrmmzBGPzstXWvQD73s40NkBifp
QORjMdzB3AHHUEUCYibXcHaTpH0LCGyuk1SjNqT3ype5xBFjnawdz/qZrzE66LgYz4tsg/d8uK9c
IcuSzGSrpqz+ZhMkT5HFob+XUiNj7/lG1gzX3EnMCOYRUgi+C8IWjW5E8ed3g1UDIo0OLq0zgmVP
WvMadSuI/v9e/HNNA1pSSKMqmPfGiHbubHM9GJ2V0YAUd/sN8xD/7crchr4rSJ2aJaM/u+ug87pP
T69q5HZ3WVTJQdUq/ActxjIGH4n8CNkALNB0/m9M2R8fBeWvSLufkAQFq/tODUqUIpcLkVnfP1n/
R1DrQan7AdtLidPJUccNYvquYwBPpk5orhPxeY7a3xE1p7I2vr4f1gzCr9xNcILVK5gGsRazfIlI
16AU+/qs2s8pWwtoHFbeaYdphVMEpqOZfxwgnvO9FEOtBp3YR/7VrL27owqavuCSyIDG5kldDF41
YZqbm7Get7Hyio8XXfJEdE+0ZgbC55RAZRXVMVfQHGEvsNunmHhL4jVVXwbiLLmisX2s96iE0raZ
CJqv/4IUK6gVa610WSDf1+VBzEs1krgPeljb64IqTbeDr72WQQMICQBQbbE5n/HNcBZJD6yXjNif
dajA7+4UCFdIAYHkG4Kfg+HDss6xQGEX5DUfuVAarcP1CJgcVSOhCwDRIQqbCNSS2biCbEwLCAjg
zPNUaEsa3zUNaVw/5SpxKSIJfOBQ6lJkKTDP9yx1Xtr1JeAZYw2/QGe/t3yjTJv9bHN++vS7PT7b
B5Hldf5QhP0kMBxUzbR8rxvIpqGw10w0M25xoPi3qowRCE3CkyAZ32em7H6AigXs3PxQvLekQxL4
UdcuT4fIkDTw88BlTj821fYyFqxknZdDamYYZ8NR8jwRu7S+xqRBVLkcRsNVpaqC+5zy1ascXopy
gXlDdlJ2jgINPy3fP/XH3+uJ2lVR/drGc5uKKxtQtgzqVuYrtglC5SkyDtacWlwpMWVpqr+nkkqw
reUCZ973/JodX2H970G4Qb9mb1qrCQO5iiwCotqr/ERZurulyEZ+t1YIeRVSjkNEoqTwnmJ1T3NP
wd/jv+R1ZbL31V3HGhlt3ztMxh+9Cdt5ps3rWhbEogwMjV9UYU1j2SadEi6pYfMNw2LIm4MD4ieD
rTTZkdeYFCouDHBfJmIz2QcatB0hON6UfWWZLUhDCYkZD3YLM2MG2Zr4G3mgtuDJ1Sn3LK0HNIGB
XZu7Ess2LZEHe7ieOqyvNwCHiqL7ZWEFx2T6p2Y/W6XDbFw3CPUNHIR06QD5SpvFST4MfVq8ijCo
gg2j3WapAyl/i+2BrVhEKic/YMenitU3Ncsu1wvVCD2WW1DUoAHmtMFxdeS6QWje1hC2BOFGPosj
+5y+rwkM8DR/77KwMAfb/XTayCML9+a2YEh3iBj3F7ZrSu6k0bD5wYXmsfUDnIhLMjitJu2oMjRj
b2X8CtQGbVd1/77HNC1I6eq2IK8yxd4Gb11pIXZEjLmoyvdfGVDgF/RtpWaM2IPRBTnGM+lMhj+M
yMIqlm15EJ3/DvZ/oXk0iWZnA01TkDBkaIX8dQnkzGpKHMXLc9D3khXM/2RZAxOcVKBYvDM6kLFQ
r+Xn+FBMb+v0hc8xYTq0MdFPv6PK15ucXl2JCFFn98pE1EDvX7BIitpOGR5tPjuUD+Z/4/1LPkmb
ZeuHBJ/MHBT8kYIA6TzJCh0KxLlF7hrJzVvuMOwTok3X57VobPvwiouMhLPln4G+R0TWu/mc31t4
8tZ6J/00/lNBUcFkQMA2IKnDX3dKIlYsPm9LZubngoH58xGU9qtPX1vQId/ec0u2VH70Bbcs6udV
T+UEU+yV7r/IUUMo4xyM1m9niHWIB8CSt5VqOlbMaRLhG+6wPMkjwVDKaxHE2IHuHWIbX0A8xBak
mVSWH36ZG0+J/r6NKz96FY6Ntl2ie60WBuVvQD9ja5vjZ2bHneXB045O0zJ3CpM0qlPvae22CvQg
36rKkiDFi9yjqIUgeYe5ODFn1HiikIWTwts+hfou9B1x6ChJNK6Qo6rYZ6qcSaMuNof65NBPY7qL
RuSPi0t49J8L0Xgb+DzwQqgItkKnm3/1hYTzF+snmffEGyQ4AFlzpE4n24MJ677g/9VD0YSOpjCa
kAgcjRZfb06QRcLSzSZXA/Vhqa3nedhuJ431j7rNwWi3C9e5Gdb9uIfI5HNj3rXwQsg5FL6BXTbd
+4fL+ZGapS02M4hGGYcLDO5/4E74ayqRGS+vn334eMFUxXfsY96sGOWk8Wg7H4m5wxFF9uujsaec
HrarOApzxPJJjGwmKGNjIHFFt4u9lNdJESadRp4nLL6mRn1k7HQ3C2mI2Z76UvbTVLmuk1qGbdqe
GZ9AVt3QryeXxSahsE9GMTDeEGhzS+zS8D2MqP5kmLS9gBiADkVEtYGUQ6miphAzxzCNMa1NyIye
sTgX0HRCcoA1TKeuRmAPJflrG3XnoMDD1fZlPfCupdzM1WKb1uU/tLr+XtVhO/polhm3o6zZ40h3
mou/hoxhI0QIucyW1tWegK/9f3fhL2hxCwcP3N+cOujBlmG9rkfuCJhUencRYNPrdwT6IXyLnPWM
PY4SK1LxC4ckvD8zzg5AyqoGJi9QpakkIEmrNFPBv+ygd9QbmcdikDlfJQu8TmW3ZW/Tq1E9PUIk
dmsuxR08DxKIwHL+XXIrBiPSM9PFCwh/amP5M4Gu/OSJognQd0X2/uDLZj1RyWwqSu1MR6PhOzjP
bqiT00a7/1DU7AG82OJPqzTaUxZkNcfjJDv9ftKPvJ8n+S/aO7Ug7tq13lXQvH00EIeDORlveLA4
5qyRQbzONSwLf1Jse8ED+iMa+7qg5Bc1FU+gQG1BXYYYjnNEPJc65qxL38zytxmvxhv2sfn4HGwU
SqEI32ePAjqLAk+n/NwW+RL7uagjScZ9paqnnPaUlg84dShjL6jqkeobo5NMDt54fxiXNBULoQK3
48Xr5i+5TLEr+ZDAe7osyf23pnxSUjYQlCZVf4JJXUV2uJUWxSRKlJjYieEAL6T/u8o9xA7meDMu
NmkEwAK1PUYLYY4tpKAE2ChLoUt4PvJ2YmxROBoUVbRqOkC/raSMCR81SsJ5ETyK03FedYGn2sl6
2lPo/qyxuWKINCws/Cc0AQFjHAhgIxLIy3+KPe/+bxe2EMpW77o1VTlH+J7relfOS8vBWgHtsHFa
bnTR7yMylrRKTXBxA3eBUuo83V3dniEZJuUBensUMbavw3JxGGBBo2RfOS62Ya4wcgONJhnf1RIK
sLG5H7Jd5IbUAN3RinAC68CBsq2xsNuTnT3Bu+kBO7/zfiW6FxYRgFOFibBDWHCBbJUrzJj7l56w
vPy1Ldu0HAPvN7lkDn/4pczce13YTq1d0S+qVimRKVrO7g73ZTh+VbNC2PpFXIoDoI2sqVhvm7IQ
kImT4Bi9H9qnGusFmC85IProqxDQQTb+uZj60QLagH4F02EYUEP+D86i3v/LDfI+fWoKD8cJXNJs
inz6tSdzShiTw8elpotgdgIUIc1mldTcbggKVixwLHp+rev+UYdf4KSH4Y/MBS4RHtFV4F+40UXE
ZTexyQ6ztSi/CndZvmvWV6MSELNOaWnyJqxJPGLcCdCFCdM9P85xCKnwB4+B7RQpLLv8lM6Ryqle
oBdpiF4N6jKJybCHv9KyCcLXeKC80UmA1ThirHkNpnAFWM7mt+FOIMIroQiC9jAi5KG5s/UnJ6Rf
EIyw49gjsBzoc38EjYxMZKvcKGmjwfPgqP/zeqqTFgAl//GB3dncLHTt2HU+3JK9kufPPQGVMU2g
WwFWIWJfiu14bccPoD9XlYI0tqKKBxdvnABkhFq++bSghii7M9yRKCqzCFqGqysajZDPZidrNOC7
pMAFGvvejlMwo3IsDwHZ5tTl5yxHWKZS1frWFKx3/bOdojbfNQhEmwdng/OKb9boufpPmTJsS455
lRd8qKSDhuyMh8/p6txUhhObE9TMyDNAQB4gP+zPrPXaaJGcn6g60snOtlL5n3mpKuxRr1Y/Px4Z
mvG9vfoaEd5nW4lF2cQRUBmnBGNmh/QQLd25+/vPM+YZtYqC5I8ZXJdEBKiZyXoQ1gl0SbP6DXzD
MxxyofaPLYozbXHZVD1JyFhcyv/XyI8vvtiY8M7Rl/Xg3YwPRb75ROnBn8taamTin4FM/sOHC86c
+SEzvleWGJSGIz2zFAPSv2jScraf2h7xLLIMXfudZr9PxZG6VmD7yDbtOixc2qAydJE/wa3osexD
e/PQyyQJfR/JyJcN6so5wOVVuCPjOX23tioRkdZW1OrFDip7ClYwIcqvfy9Yno9HVsjVTMos/JQQ
wknbEGK5q3+H1T5qtGskHaXF2LJgSyvwElC+kt2Wq/1E7m3RvgA693Mq3OFo8W22hfDVzfB+FcPC
dxmslRKMV3Hf5zQ++0uJGufrjGBFc48xXDNIr7C14bviywR6qUM8EI/1jnZt3/HW46gFj5bof4w5
bPsOnJAcSlBGVAJ8Mqv8qk/F/cE3hpjROxkVCFq4QYQWQ4lmoZuTHo5helVlCJ8CYrg3EdqBV6DH
koj3WeGzmzu//h+Kjrsi3H3YsG8kQQBkTuN/x4IacK/jY6mbwSZ7P5zDCNDm8dWb1WpcNiJFhbet
80xOLssryPUzjxLNAARqF6oVeuW/wuz2GfX+wGRFB7PTAEwMnKDkAOYAt2NTJmYfTnN8Y4LZTEFO
o2mHxx0G6h6WFRDyJXWxMXjNdhiW17ktAk/n5xW51T1ej7f2pQ1E4mCUPR6LO9Pn2LUkLkvMuJ9D
tgo604MF6MK66l+NqEcjxmU53ZSs8MkbWjjASRFKmEHkRafeuPKrsh+K0sOt9OCi58kxwedAg8sW
xctA8ZSiDdEZxuiKjn/99zEwuy3/P4E+tynkTMgIcQb1Az3GxwVBRTrE4vDZHZcIFsTeV8xjK3ub
BMqRgiL3JURGmPcDpWfuvIjtP2wbnh0R/jJ8VRb/k/sPgKXg9EZ6gC4XH/XWDBbpDvM7Tce+X2Ng
MCpvlcNfys2bZXAyNQr1ejyW8AHCC66FqQpklPbNgNlkn4veTRVjMCI/zl3RTndshiBYo+nPN9go
zVoOhoa/FQGJzcF299kOjvmq6cNmdfK6QHOyVS56dsna/ll8Fsp1cZG9J+3Iy1g1/83rwrOVOYz4
ya7DyEL5T0kagY6sYOKrjifIxsWmQz8JwFV5RgC3nn+GcqjwKsSFu2HUQk8ey8uNJ6e/psj9+BXt
Wz/emHyFnD+CHzMqPmS0kc6yRrpm+iMqfXR6EVf9rqIDHXasjiR1oVspnm6w+cjxvfTcahyxGhB5
vFv/LgpXH2fRQn+GZFPYRKLxMAxBs7Y2rE10mIJvk9cQM38z+OMijbZ/ZhI8hJj6oJpcaHSsEtxJ
AMS88WpzALnk3dHEkEZxUl57S67aV9Xtkut97Lk+5fUq+kFI8d82bXI1RmjAH4KNwq7XErbx0pli
obB0Ru/R0rvnWMsjjRznXNCGeULguptWDGsvXV/tPYGcgVG7e4cUsgnX0qQlDJEVn+vhQAcjrCTf
k2a8HhkZ2xUsuY6frWwNmRIXLD86/dQ3mQxrZT/H1EIiVlC8mvGXt5MO3lovGZULYeSgIBCai/m+
m5DXYcrfQAE4IKtsbGVhMgrzR049MjbTESQ+z4L/PZnqGzzUe4dZbIZCf+Y3hVCcm94QQGA7xHJD
Y2AIa3Fpx+OJu5r7zGxsVq5PjZPntKAA9akLOiFjm2CrTooJ3evT6GTFVBABuRTWobA0qinmX2+F
8Kb1TlbbBW3rxNtnhlofN62AbYVDnCNiJ9tMTqIKVV6peAEH+cv+S4pnIGvQjE9lMOMz2EHpoFhr
7gfItYWJXSKuPx90jdZia+yZLezlCywc7keB2Jxpkhu0cOCHFpwEZIZmLEJzIvH1DYJj38EOn3+r
9mZ5Tc6JcMjiKRWhmRysdsj8MbfRncfwXycC5+vTqKUHzFUwDJLbZZ594UqRdNqdVCJDltYt6xoM
6Yw1ahKDXxf2RS588srhcslfvj9HT4BWTq63+bTl6XoQorijJ7IKcObXFstnXMs2icVDKrlrctms
a0qKJNgzkxhwH+OczQSeLTSLojqPdzTNFGLk0SmYUKTJ37R7SX4ruEp48PDagZ6R7s+LQiX48sJr
vsFcB8VXjZ722FpH3Dhilf2NVyFuR/B5SPyj5Eb33k+7pR6JdTsVcwHwoIFjf4mbQSZSc324iYXV
fgBvFFIl/FCI0k/czLdOckrAB2oHA6DeSXqFX9ahDENXelewrD5v8opfJhQnu8Kf1Go5GwNcsz2X
G8DkXVUuovDebYgzD9dv/sZmGWWvl81EB2yYrxxbAl3xKtiG847NA+ilOiX463mr99U+p1RbFUe7
X/6h23FxUj4ztfVv8j0ZAT0zcO7ns/4zXzg4FUwTsTBW7g84mAVw0JBDwLaL8cY60PLCh6v4dMbm
mspOT7DcLBOk3wXi3QXrcPrqlSwE3nXHx/TdylhDnXi3FlXlpFLOHUXezxPBLT1uVAZp312ODjE0
n6t3c37sjFJdnJcsK25L0/Ih07GUzL05vFboZreiBeDgdy1iZ2FRq0XqLhg85T1qJ611eh2DgOYj
op097leO7uQ1orDeXgtBBltI9D8pCbrnDrDVqfPjy9hq8TL2oAK5I4J2gUnxP8QiJmDYGodpyzOW
jLHYWS4/RXsguY9EG+vDsvLVoFbs95iso5BF9G1YZ9ykn1sP1GNlBZvMqCo6sOpgvfCEGA/OkRwl
6t+YsKZGORwe9j3bsnpWgc3oHF/z/wyLH+UnGgRQKEZRaegjGqqZKh6yAahiqsknDe1R5OUsOYvZ
XC4Rx9/dJg8lnDTkkopOgNKyGI8F7k2CYy69XR8j3NKWx3RI9oS6Qwevzq+NzR5P8Zk8hXNKV4f2
lWR7PWHJiqODwzNm2GttBwWs8S6okdVZS5xi6fbbpmOSi2/CTybBnPVv9BDPWg9SWTUvwg+hLUEb
zz+WlrEUVTOKA+vxJQKgvS5MKAS/uebGnw9HRllIfoPfuwG7UgoOAX4NGwvu9e0MRrpVMFHHWECu
JzPBDsMI5P2efMovcFHhcipoUFc/B8vX95muQ1dRNRRwH8b/MCF4+zrGK3IBHFVHtHZ0JyJVbLV2
XBAHpJAQoqALsJBCIjG2VX1IWfth9usugnp0EJtOSASwUvaC8XJmnRCa21rig0w93sYfOqYvDbu0
FHbCmyuNHGIotS4iqESv2ZAGiVgNkgAiNq+mBHEdJzCBHgnN1arsbz8vwbd9j4ymbE9sGQOqpl3j
9H7cHBrvFGrtsbzv8WlMV0hqyf8SlFEPvaqh1hDxv+FhhX+Q9Xn0X2lQFJ68/uvn6JHbpAuPC6LS
BhLHVawvKul7IxC5sL/zJaN9ULHKdWkNFMm/ulaQB5hmE14qkbp0JO9ja3Ry2elP8sBE0lezpgU7
oVCXT7C0il4ngBB/UpOCB3c892S0D/W8wHOkBobeVE3W00X4J8YiGfy/w1i1i2qM5fZBkLd/OMVG
XzM7KuQ3F3fAl/DK4JgcKEYRHZcuyA5YadweJ7DyMonyB8egWS79S0cfPRc3tTI40h1De7Tm07l1
qBdJ740Wz0u9qUgBoK8H0qS02LD0YZyfP+pp0sg//1iBC/Df6RezEWr5jWDIpXqt8FJV4ujm4bI3
iqPkkJa7olsJv9F3Kd9Hm5MPamSlBwAXF5YAHW0JH8eY+Nd8Vm8+XKj1JZsGsUAOhii+i7TVbRbn
kxWO2krPVzspnIruUZGK/4SD/W5uhsj929CNRue6v9IGLivGEIG51XfZ45G2vz2eWEVQfDBeOJoF
ial/HipS96tI3s75jEbHxWLGb/Md953u0D45L11tusinwdyjXo9ucu3S7L/BNLhpX1QkBh8zk2br
Gq399GJYqkO8eVJwctPvi2YP2ose/z5ADMazDbmqSSm6kb1hI4UaaKrPHTVulMLJgjpxMXAnwGDt
ePiIs/TIGVBWvquHxMP4aVB33xmefDu+/YUbaXDrhJmN05Nz69PCMTdeF9panz0dTwmVPbz6jjRx
D0tVoNii5PPRy7/V5FO7NhrLk5vmhpfZ7QY0PI2JcAWEl5ydr5NrlKp1+8lBrMCYoz5Edjz+Wf0X
BGTVyGJLxctMgqQc1PwTso1lFfDR7pvKoJN0RyAWAnivYUxtpyMqryM+XQ7GgQGTRkILTtjyFV5U
kNNglFkZgk6eq/Lin9unObS3cWbD3cX0MZhXYcNonspvdOsr7dm1O0sHcaNzd6HYA9zEwOI3UaoR
Qkjzbzr/+3YZwbi4/ZAERPqngqefjzO+NsWV3MMJorDaOIUYAfHvlBoSPUi4Ix+qncdg9Hy3KzTn
L/Ed47FpbA2VZ8t96Kp+xaQZ55IJwnKpVokzeRKs+yEiJnOZj3xwMOFfvda2+3lx7kEUq9CsNNcr
0u/ueKivFJWradHbFJ2Vzz3vFGS8GcLeq/AKMsGqBZYMSerJoDXBSRXoGN5mtBCgiq0L4gpWODzD
+BB8yNh0oDK5J2DZ0BWkZqJJd3n9OCElPC9PEUWnIFSe5ucf5wqxFHgCGQ0WvjVzTXTl2PVZjfvW
jvWgqb5Rjx9WsvKvTDve9QAF1znpLhPX9kyISCsPrEkke9KBKYPXsnFPhsj3+okvAahiRwurr26V
vL7xoBu1QeH1UAYZVQBp5YSzJtk58qXCUV5NhGMdsvNXYBUssDaiJi35Wp8bjRgRncKhLpLO66zZ
66jHVt7HLgJQmJDALwoHpROAp8C2j2kTChj1amflfSbLFpFf4LFbYZwm0XLw1pj1oV+YqVC96lLO
BQ/wCxFj9G1eWCMFgU+sJXmAg3Jl08eLFUUB2cvdcwP8WoKfECllx1007zQjtHQtQG2tPTdLpYMs
nIXIPL+OfOpCozyIR57hZFMR7/O1gRAVxBg7I2uN+Z72Fuo39uCAFXhNDcUUhGf5UmY68UFHiVNj
fw8wuofSPg1a4hk/nqsKpzDjEi3biSXtGNvXJ3HYuNazHOzSycWDCTEbFvsXxZMSfAZSwUGvFkIH
2oh5qW1C+pianKNRxa1Y106Voipw0WghGSlbtXFIBxt90bnYcX3lz4vEQSpoQvD4ViyuiBq8JBDY
ftSZT8HQaQjYU3HOjf5owthL6TvdTWeS1nCDgdRT6mpo8pTd9v9v4JUzvq++Nkp+WOJc7E4m6PCb
iINy3enHezBUyQ5Qc5zllBvdeS6ZgDtmTHmZVPqaT5yyZh6EPL0oI6mEKQN5riA7oxmSBb5BfvUf
s7U4Kf6ttjT6dOn+1gJ+AXSL6oi3tjrPMLN+qdpvaNpdyIOShSXJrCX5T7laDGT6kAvK30FiwhzK
sGIxilu+zkkkov9keyrn7IlXGP60Gtr2J0xAcO67IFuN9154kU+17GoVLSf9sPNM67V/cN1ZFuPM
MLhejsFE9IeZ0KBlQQDSYhJPmi6Fby3oiE1eQXAs7umQVr6E6/uEP24ttqysIKooa2tFxQ7W7HMq
Tt9p6pfDF6rfQJqVpqbgHyQMH5B9+0YQ0gxNYDNn3nuK5xdTFhiYEEWG0DI3vpEAqN5aCIxR2MiV
y2RTmNgP66FX1HiPMqFLb5BhLwcDqqy72TVP6ZHf8ZBNxkLjahxkSZSjqydvYfinef4eNPc73yRT
X79A4cAxHZ8UGPcInFoPgHz7KULe8B8YD8GWS3YQzk1vJ9tdfcKe/laTcFb6zdXsBhRqL5lrckpm
ze/LR7tMrvEfpUzss57X2DpZALOApjq7C/oQciZfY/oiJdD8i+1x5g1i40IQu1JfOf5HCFfTzf2R
YydS8tGFWFkgjb4FECCrdmuteyrGZsp2M6QDZ5IDaqZX+cqnVQvx9SVh5hRqPhFmIIKgvbKWDJgq
TPuEcrGGFimmVuc5sMbSCnRWyYMksEjPjDpeoMAoWDj9G2zVdtl2NN0OTJw6/XjkQ0Isw9m1qKSn
S+nMpYAUS0GzHAgIbHIEyQkiN+V522klnC1+2nmZYi+GLue2my/OBDMurg+YXcnhkL6TUg86LLr0
Q7x8SY8WOyVYqhjczV0EJ+b4nB0OJZkj1khTq/NIt1++njWmGNFBBwseUHm5Q2yt5YBlDQ6tWn5G
0+3WTo//iH1lAXAaIkzNMUX7NCSC50UTiAEr4Nycm3a6rFSHUCFYAxRkGV4kKUF7M3SH3Dl44mg+
71A6/qv68CTjBA+bBTokv4ndtF3KTtvNm14zVT7lpyn1pvjoIZHsTudDTmx8aNVWvluiuR3ZhCZe
bhN6iRssj+SaK9FzE6JHula3/yHywuFG+MUZy4MoRJnUDjPb8IxfawiCtkfHcLBDNtTii2bglVix
JS5JoAZOquTFAMTfEQDf0wSyEietTcTF9L0IHTlx2X0H3VHu8BO+aMaTALdmTKGMh/QWO1Zenl2p
edmxgOZiXnRHdFRNRorEsu1Qpjw7MJCSQnSqm37rNRjh1KyAasLb7nY+Pk8vSyIsLVNzHcpvH1H6
TlPkeD56Hv/6OjoPd/PMR0X/UmyabAr+wwd2NnqwjMmI59BODGu6jw36GCH9oxrTjI/LkU1DzKEb
dt/L+ZAiJAQUnyYz0NA3qgkGFf5+POEvx4wIiMxikxaEDgdkutud0MInO++J2IyGPt5Vqed+mzBf
62psP330vT6bZ1C7iSQbUYZm4whg7nw8hd0DMSg8Am/9pMIhvDZwNZuM7wkkQAjWKV6cx72lag2n
I7bUPemZOe7m09LiVuqwacCDhHPvFjIzjUfyzxigWnb2BGFkTTwEjfvXnBZ6r2Zahl6neI3ldhfa
0/jlIzUXSooEgmz2m10xSyzPboJf3OUx659HI0AIgQH3fGp4enCkfer03OFzwTBbma3Jba0QS8Ip
9Uj591OFHWrQ4W+GuFJDjPgO3NiW+CvyE3d82rDK8weDp8uD9wgVglGXsNXhyHCBCtPyuQ1yFnH4
I7N3YNOoM84RTMqhmI82i3hcsVDGY0Bg4SPhzyi5G1Q+VfRtM+ECtVXfVeB0qNeQCeoUtxgWqLmb
dcJENWZqFrEyFm3ObtskjYpgMHuqxe0pdMRP8pks/UA19KsK3rsffqQ9UwFO9iCsUUvfODcHNxc5
KNhzeqd+N1z6EvsloQ/S2MSbhEt9GCEGNURfPYYUalulDjmWAm8uOQnsCqqSdHQAkg7/EguTma0V
AuFpOUgYRlvxg+qjxZe1SnTFAh8ZMVB6tJ2+t2+OZfCMwLOmnnG39/hrPE1DVxgZ/us3kylSeBuu
k8OFj8kwn/FIW/pXTAmXfsoTWJOFcC8g4Di6l96AqCB9NpJgM/q9QJ6Ns/whFUJjvoHej8bJg+kj
6Wl0A++pc4iO+Ne5h+slj9Sc/7zTybCFMF/R6RF9XjzjCuLnG3ja48+hDwdTAvabOD7G8h2yIdKW
g/1xvC9cFzRKzAFOyYfT5eht8k+bVm7IwngM+aG57rLq215E2ar1Ozs71EXC5Eq74sPY98mcxsyf
324yHvvOOF05Y5wK4SHjrhyG3panpq/Kh+5OvkIfB7ab9y4Bkaj4nBH+WD7UrV77YpLyWKLXoHC6
7NM15+ToLws3mN3A8o57MFPXuOaO4Iq6AlB0aKKHA5NSn+YJ5He+2AljeP2WBh0DXvVtOMMuC2Zg
LUayM2cGr8JJQgr61Ozx8J2ofBZX6gipFZUnIVp2ZSVTbJfWfXGi1W3zCIRi8ByO7Exu5tS3t1ow
2qJzdk2coW/lDKWH4KYQ3RrEN2U025h3PU3bi/GeKmBUgdkZK4b7LYW0DO5LoQ9/U4aThbHNdYNc
yMjggXqPwL7Rl/D6SbCsGI9202/1EvVSTIgTa+pl1rfpxBy9A02ZLS3VEXTgm7X1/29wC9deuXYl
ZxRdLZ793W4yN0MdWkOli1aCsq1J/5Y8W4xWXQecGTxwhroucTXS0bFpBL/TlFCV2M8y3BCrXojy
LrAhIn6m0zb++4TYRyQdbwA5K/QVtSYgjYi25PbjhLUUsV74x2iwOUo77dK/WQyf2sPYM2CZmieb
RtJApgK8VaTCWNCtWijpme0/40vwxHkGJRLGPB+NHvy+jL1o83EY59ZRoUTMm2ADh3fM77Xl212p
1wzNUUwH9podkVHN96l7h+ZQ9+wsVKTpeM4sgqMl/HU7wrgd2RFr1+roo2v5bsoNKA6Z+1V+bPBi
ryP3CxG1wd0qFy1sZ9YuVsq4bmWh36f2RII2OVoFIyplnEqNjMFJzkrp8UCymljV2c1wdhiv6bRe
8a58yIX+U6h13i3eG5Q/RpVGiIWYwwwtOJZQcqmpKIEULxOJBJS97bRaUZnVMMZ+Caa1eespSotW
s3bH/CGHadZTSQu+AthM/3ZAvVEGEDnO/DMTIqVUStzmJJPQfqhOrU3mWl3EHLC5YUaUboO0Ypxw
hb+8lzXig4iTpgp1jqhE8sHdaMCnnMTt4kFJ59DmkMtmvMFfozXkal1f8f13EFw4dIYz9SyHcxHg
BvQM4+sp2vsVlhc3TnllGCv97xt0BDZEP02nM2a5bAUQa7rE+MmiITMThAULY5O+VW+I+FXOVYgK
ixzoQifn7cPrCy/eY6wunRS/HVHCvWmc3MX+deWy3jZRmN+cNuURYMYSN75I3+Vsu65WyLt+E4TY
YnaUMZoJaZJXoc7GOsz14rHiWaE4qGM2ycJEMOW1eyWKNKxIoertQw9XWZiaa61Ktns4JVO9mQRA
PaO+ReCDLVCg9qKGPwXr7KTOnYvN/5MUKxix+apm+n6Eueu4lZvBC3fafwA2InvcHYnpPUv+V41Z
Es5dqk2T529CkTfdyzYLy1spWDYsBR3sbdT9Fcgzgnh+ZO5VP1oD1UB86v+0wVxJ5U3la/lo50WN
I0d4Z9dF/sj7WRP/g6I4MQV6hfvPsQV/PFrBWf/AIkP1kZ0DXyEiP8WOO1UFEOmKXDXtjne40K+m
0XlruORdms2AijyiwZXTEa5wiSw6gzRm2aLiA81MSh5iNxOw7xJ7TFKWoTwqz7Gj2YQIdRrZwXgh
iQ1rNUv3KLy0eclSaz7Y3LIdz9mYPs2Q0NcJUtofARZq/GwxP3Zx8CXQzGvdySqJnmVfstw01CUt
7ANmrwnPgC1rDEMyxD3hVl7INEVc6ncfFvssLDqPpPd5m3ORwyy9PQ9zGMCV5mPD55a4xZf50Vsj
AmOdeQIX5wCkv/UJtfbJjGLBzXgOcDUVSTWNOnjwOWtuvCfSpoEZxY2AHK2qJnjO+7d+RnyYiz5q
y2143aJL70V95y/rX59GBsCuRl57BKzWfx3zYPpGzOa+rF9gGyWzV8aLYsAz39WPntDJr8jyZQ5n
H31Z0Kqr+SLI7suW8uSgxdu7sS2/ey77oqHCpD55HmbZHjOsHOmr7Ghquhdp2ugoC15loQmxcCrC
kPr2Ziz6RqRvvFA8T2GWacuiGZae5oxYN4DwDYc7PYBa70Zbb3JV1b55mAnpxYIPBj3Xx2pBkSTE
lrNIxDyM1BU8vNASaYqLol4JqYTa/oJbU4uJ6PNxANdg9wQk7fUthBQJj0QSJicRCJhU10tqk0Ue
bMxSS19T2t0ve7WKkO9lJKk+m0ZU5Q5VTZbir0gox5eUg+dZjJfqB++6DtQVV/cWrCLCSoU7McpA
snCbdZc/lpehBywUkF2YtC/7enFghdTe/JEkEvMmi7ZFzjT9M0eOi38KQWJh+Q6BBgLOMAvqvbVu
lnpl92SzKTKC9NCOExTE1fW/ZiD23CHhr9qEEsdFamyCA2CAb3ny6vFomCsEo1UtHt+D290N/28R
tvh9+xe+Lz1bZFDIzQVYa/iBa1po6QxzS5sBbwSInQ9grHf8AoVsz2ZS9c9qtT+VKTc5KRnG6ZzU
9AbaSXhjPro81Wk/13h9Wl9GQjQFdnMJGbXtNWZA5sLnvHRivIzIwfKSOxBYUq32hsUp/tsnTxUX
wakysMW1KLbZPcplZpqcIE7141ywp2k4EbexkuXja+gT02VxX43dydLqPTJslQz+eTVgwkHxvQ7t
4pS1Ka8CNB2BFUVglIXmW/S6AS6+nDdtpAwDWEPVvGeIEmOD6opGuOL8R2zbGBK2m7TIx9Giev7p
W8lRV19TMcMxbV1A5yJouDsqP/1+1VMinWNhA5W5vjeupIWnmPUg/dZDZPeIy11RNY8ZiTKRrVDA
ion5dyjqkSbBuHYNf76aT8wTpM9sLDC4c8u8ybvXgs1g5tILatZbGTY7amZcivAdLUQA7wKIJqZA
3qZ3PN4nbJkBRgSVw43d15p5iDnNGCOWjIn2erXnvdY52xSBbFe/IBFvw0WgMSp+A+HM5+u1nVkJ
dp5+AadIgQL/dJb0F54bTBwBcSYsRfDWkpiFg4dfpJ9cC0KKgW9ab8YBj3UFTVdPqvYW07Pnf7eh
hD/Uc3LYGAPDkYSz5OdKgWviImX7uzLyQv89DrWQsbZhP8XGCBTPhpW9yM7XfFCJw2pWsHBVoSjV
wRt6BMGFolJULyJ97cX6gnJ4PLo4vMcLDLRaU2xcDMlLGg9vj0k9Sk5wIZCsTzl+zcZiISVwgUnm
90BJPoW8HJBHogDkKEHosZ7o+VX316N7SR7Lb/Xx9cJnMwTbVn+EON/DNdhcqtXFwz/Yf6ACaNOg
fd/q1DYjp9wA3kje049ma+8q9ExBTGKqtMoOL32da4MPl0KhEP05nUopt6gLLVAj7vWjYX/zZmDT
smpXCXzf92U5CxfPhLw//jzQ5EOx+yV3l11XST42PjdgehG004/14V7JlKtoOiM0XCQaNqtlnOkP
VKnc3JsMb/0U8C1u7O9//6yHLwBtbRnBiRbFfayfC72UnRPQl9xcFZcziNQjlDc7jXNetXEEqpu+
QhY5wFWxakwDOfQWmmG3AfAV8JffYSBipb9Gz6joHqJJ4T6nSjem766o3OkkR4MTKVJM034x9L3B
Ari6pC5s+pEV+hlUC2stE876vdbE9pFGS4ZhrW/IzeKXAt32/9gc8fH2nKjzFq5vlDXsXIZpRp+J
mPMO0nXrm+8yMRHmXJ2O3RinSCeD/oreC2iJnJhHsWGUOjNjNVL7WFDZvGa/lFrp1ggXklusujEs
CFXkSf0R8JnufprsQATHJLEbHIv5CU1FjqR6z1/48q3XuU6+1/rPYgOjSxNIw2mZalRvAPkKg8fX
vhA+ngwjsqdpSzSlOiI43aD9ZqapkvrdBf4f5+/J8fljGDPsDHHoo2bRhq7V2GOJMZDBHGuvSSID
L/4k9XiOMFaK0kH/59UgBpMabBTd9X4TcNJRl2zI7SgwYQYEJkBVzli62LaoPDYcPKDFBo7rL/QJ
qvoaNXJh8ywVHHOu6TJz+U8nrYg2Ce6oLwA4muBO209VvcWGHTV5Srz4QGDhAx6gEhSN9UpDaYHJ
Cto4cOprfI9Qe7fbAbwBXXkpjSBaRbkX7Yi/PZ1qa16NVKSg3fqyDyP8592FGJZPwU15vHur5vHv
qsMyyOki19ZSRRWAL+H5aqJqzyYT6ydmjH+5yBmtDM4sJHa1RFjCNV/dzN0lNBGXYkLrVJ1WeBHM
I3S/JcTiHcm7lojONNodxqFQttKRSMyOLPlNjDZXdE/a69ulipsHFBaabLjNpoq2Unv9mJXM6vRr
GSKlCvQutoVFcDiNJSwY+o2JDV6wbFG4FXgV7/8zHmTU0vuIL99aVYrNdSs0bbYtWQa2LpwhcySK
7S85THqEzaoFCWruNQCXWeDUtO30yu5g81UgkZTgsBAvozKtWotzBDIgCKrroKtPQwKVd/pwpero
pMLbf1dEXQeQ8+ib8VUsmR+kXYN7nHnetbYGjE+sONz4f/2vF1xfeZ7LMNGY/o9wujaZIb3+Jf93
mYVdHbgHIAgSvBb/0pSYmBPNF8nkSAwUyjUnG1kX7dQnIKldOmSuvypsvDtmqs+cNGlZmV2Pzq5J
nXr+xUIBRn+u5xcbgWaZnu+Dkf0QML0TSCrjtDuVyRSQ3M0eUtmcDaV3C9zOAt4OzT0u9LI0Ztxc
wfUugEG1725F8/Utl7hCw+PWi4LXboKOSWtxOgED93kZUn0jn+Unpi9P0b0+Df9dPgXFMyVIS/If
71s0MFSUbk3VHV+zQF7g5YeunmE4jrkFfnTmLBnpzgjqex5Jfc0JlY22CcmJSxbHdFYT/5zBlWxk
55NEj0836HjTt8bEBqkhFfO2/aCN6O5AlqDN5UIDw5KeoOrWTlwXv6f0hVUdNjsLgvqY2AiIKoNu
pBH9CdQcqGlf0Cda+PS3+jrg3blqZ5ERsyInsvC4w5PozxhfpOsRNtWm2IlmLrX80tQxwWu+/0oa
ef0L+fM/7sT4LBxLqAr7sTCcJUgxM/p8E5sk6AT8j6gIkcr/D7WugIcVOdUzkM+FXnNldD4Bn3Db
0aOufP7djEDZDZwCEf3bdPQONhTRY7nGocl3u/BWG1EL6kZv0w5SsFgrCn2L8ETTsPHod0JfbTMI
KtL8ETiEuaIFpo0cMbGyCZVJ0HRIsloi/htgfUY4g2dpAUlNRXltGqjYacnhKFG6mpynxCn1kU3g
VdNQNSnrZoETQ5VkowzLZk8kpte6HOfsXbyb4hRPtdQsZgnWqwjHlgJG3xzfanPUTqCSGoCr0a9n
EWDRNwS9z/ravmLwEL/clUgYHets1fQg/ZaZX0+MnWyerWbx7Y3rOG8qh4VnknIiBeNqfbKgeOsR
0BSfrnffQvqlTn+YJl9LSe8Ckj0YzLGUIaHTdc3tuhkzosZzUgG3I293WDdfK09aQ7bNe+XDfyAW
nJfx33QdHSDanzmxDGWqS/R1KkgyZ80gAmQKrriWUCcFAZlArQ3nfcSQ7ghbMwFv8rQ94BFFZcGQ
ovUGawEywa1WYTCuvGbvyREFukWWFa6TpJeEPKmaomBqga+/hzOc7DzF10bGGKtqXLFK+E8eG08o
q5LWYf49SsCPOWiJXIcZP4qyRSg0yhRLydnDd9jSwFmgqODhutYmYqODwP3iJZJl1Hv5rIXuZpHZ
85l/O5xYBuDikcH6sxf7Wuv7PhEbv/eHmoTbieKZE/7MM0ilLsNWnsAA3uD/KgSnk5uYiT8A3Xu9
dfhZlB7oxdNSgY2Jj1dCyy4IMyFD/tWJXZppF/QZkaPvjVvkjPn/rR47CPkRkZ+wRRzDuEHrTDhu
6vdlRi9UsyUcF9rWh5LQ+uP1Yfxq1UlJpBIYsMql+3nyJLPuA7VuJhqyDvAZDQJ1htnxu1n++zMJ
YxC7HQbCCqW09SS1EEdQmb/vb3tlD9Yh6mBT/mpLd8OrCJLhY5EsylC2R84Jlxf24ZnEJyy65j9h
O5ItweOa3iy+foIL640MPfhFq7hhBDSI09jinf/XdBErYCONCqbYQprTjWUPhwSxqA1knBx7nqMa
vsWyn7qP1UIcidPyMwc8cHUYuaXLSDWF3GUk1dw8sw0zx6VM7DwiYFu/3VokASpgAbX7qxeIsNWK
O1f+xqeB+l1Mze0RZMDeI7gq5arjonP+Xc28k3V62XznoW6xs/MaMJxccr4EgX7pwNI3Xb0dV+zu
XpP4SG6KHp0R6DBFKn7TzBVcg5IFS9t99xcmR8I96Oiz7IM3FdG4F0WmJjqEJdyRIYJIv/LvLJgC
ArRRiZsbKyGRK51JBCBnEvsXqEiugglaKwX85QDfzsLcAFeb7fb8KVMhkF04e+6S8P0cUHnFug0K
6wGFfrSRiNYI762MsdIDWtnfS/Wv3YFILUwoL6sORhRvxPeWHHFBYhBxm0xW1oxdAwopCn5/2YXT
zerzB7OmB6FblgUNMZ4b9EdCtVxbfBUUWjVQXdHrpRX37oj+eUA/fglOFg2r+LbWYeUAvGE44ClE
kBMyUln84SnS78ssHSA9oKlUPNl489x0qfE8DPetPFyFspK1oKevds4ub3E1m5q+0iQ1uvxTbuZp
YdQmfRInIT0bGb+Y49fnsLtyJxTC20nBJ2vMFWzNMMJXw9AUPgQnzkKP8xrtqxdi4E9sc5FO1+Xj
E3i6zpLiLMGGAsWUs2EfJsYJn6ZULSuEdjNoshukLKqEYGf2IwkPuDUXgKBWsFQisI99ptEFVNbV
0/CNpjnQddUF0ltWfevjySjVuN0WDT3euFjLCtgGHmq7+Jl0jivftlaA2wT1f0sIvuyHI+xXid5R
iziDulL3j/FDhdQVp3VAmVcYFUMtEt7fiIX5pItyKRr0IZSp08xE1WI4hTbo6z+XyBW1fIR6863v
vcvh2cktO8oPQ3K8ioIvR1T5aMT5JDSAp/9fmgehgKIyXD2TNtzq440zBZtnP+VRY6wxHkLyxMkX
qebkjvRQBiEmRxpOoenVwsikZ/z2QZmhP3OrYbtUEtbHGgMtRHYglUak2KFQP8lfidfVHWFyXWeH
Ol4uLHNJXJu9uCZ+MGwTkXLye8/PStvpWR2+rK0A+ZqMFCItOSaZRehH8bQXdYHX35v23d89MxFG
AzJj+cTV3pIFW5S0dkbUvmbJc8m67zmI7PwCDindglQok1AqHjEhrAV1VWb0VdTpTGkHv9ZRwjMO
J8AvD8oB22r9fIMRqWFxCQhE3BhueWbOD8GLIDwvr1C/B09KKuiWOxtOjOhvmLu2bhbu8j15Q6g2
yJ9Bzbl6HbpFXhyIUq/HHs7ZR0sWWHn5RNcC1FcljF/D9l9VQfYTPWpCaVTwS3We7vmivbjdLYph
0NxS1ygzbBwSLbd/Xjih22jFkdEVF2lDRaUsHOfi5UKB94/ySiSMjGCbsiiBytyzlHJs7RpxlByZ
nq+tdJQoEq5bc4ngQBT0P5+4B0LtLdQuGhk67epDWpz54dtBV2d1H90FcIA83RAA956HfJUhwRF7
R2sqjFoR988zxDKH5sbQnOGxEa+jvvygqPwZFZxBQ35CLqvtkfjkn7crEs0Eu4gD2LVkyQlOCeOB
j+hLESAl0023hhoSYWMgGya2Got3NnCaSkUYYfpDQJM4/MnCoedzf777mu0Q+DzDn3gp/7HlEE/D
ZzztW+wvV9rDdNrfMIpd/yi9rg3DWGQZ5wcZPHV8KeoymCoNwUtFtUPiyf0ZZ13rfzJnE23+5YkB
kSf5Ldc+HVtXajFbUgeAeq2tIWLmYTM4LCD5wIV5AMY1nayQVLi9BcW4cXNT8MRYtvcQWRC7qUsE
GeHa+xehtnZklJb3c6ePfTsmlt1sgNqllMGBMmjskj4+GugewC5yrTdHf2WBUDrchv8dB/nXMMX7
lY69t17pmCDJ1UEDfb6iOCtgNt8qlVZwYotlnNCa8+Db9H6BihNgxwA+8JszfWEKhRScrZsOlQr8
9MP/23oBKEb/2CZ6/gfREH7uYxDAv6WB6yPAwPMP93CeFuBjhLd49B7CSsHhPK5yk24Eo474HwPc
9R9yaDTT2QXwOuQKlytzqJjQ3VhvNh0pZtccwo/ZB3RGi1oRu+tfQXO9WUT2skOYpGj4HqqOWjga
/eq80R5dlz0IhO+J0f+l2GMPJBssplZCYMTNaJhWqarlUknK3optAkb+2jYsWL97C0cOfOH8zJ47
zkbpSA6AHkVdb5xirIwMd5XsumZ6yb4+/oznVxLeN6PLrmS/Ed3Eb5kay0NLkdJ/WA6IkkMvrGiO
6ZgSe/GMX1j1EDyDgr6du34QW8Xc9Q6H7KVPsqcQU0ALbY0Honw1fSRH05FBPV5ukoIJOt90+Rj9
xH3H1Umgn5kGvD1qJnSd8N2vkg5uX+pNbYLrBGUQG7/JMzM++OSwSohZLYs1Yxhz8shoEPuH/V5T
PZagYoBNlHyxoX9/Qo5NVzEiy+JVyWXpQoFPHvSIJtPPi8Mdgk13950DFebxyxexDtX7ni34mpj4
G6+hGOK4K0ZJNqGNqTc/3ksfH7GTLPbbrnHjpcAKHJPJjRiU9WXL7ZLS33CQBSe7zFUby9ypraf+
QuG8mwZ/K0mYhMt7PO6C82QqtWBhi6mAUdtbzKeMNh+cSVCdaMtATJ+Tkyz6NtSe5VZKX8dOD8El
7rBix8/0UOpq2mz8xM0375hmibncKYwziaZns243xTRe9/MNwE7ylFgiaLmCXZYhOKoG/qwzvwVl
5erBhzbO8bhAEaQNv/KG1hfwLggy32PI1wO5XXaPnOTqo/RJKeHdaEQZjiwjmJxszrZHRrunkXJv
AgjPLSrGOjkWWiCyvLY/MmCkFS+gxFvRdjVIeI5OXsRdtx09MI979v5EOy/kzRyPQLLbwUQS0YM7
/T+tGaS2Q5NHqatkPk68WiI/y0oFpUabh8/R/dxVV0JsL5xbdHALwqmAYqNIglyVclAj+SXYO9RC
7fmEdjssfM0bPeg2yFkTEOSLmIJ2/g4SsjNrk5qgL4VexUGlo/yAq2Vf/3JI6jpgCNmW4oAIX/u0
6+mWVviRW1tl+mSID4LuvIlPN84/UGdwsx4s0eR2pkdDlX3gDO0lEK5R8YbYycLtb1ioV9aA0lF2
hl3VcfFoOKDFQarDLDdARPpr1aKaqj/TQiPCSVMCKLKpm0UnSrrBbnQ8iQDM5VvJY61M8QGoOVB5
3k7vI2UVGdZOfHyXFWmSLSi2GRWgbnrIc4JlIxDK+yAdbCb8bkxz39jjCVndsYpyutAAHL0iugoT
e4fjkiRiXlbhgY1VO519CAIGF7tToFPkMk4vycK1XSIC/gts8Pb2XJ5Wqw8ViSQwoXwDD6BR6QUf
Oa+1pS28xpTF16nHiDFD2/P8cIMYQZ2AIYf4IRG2NztlNdQqP3wpsC3RZNyAFOOPbt2RV6AZKcdW
MCzAU0EaB+0RVpm7LatxVaDP23hr+9PXGUrY/1j3aO4PSr65+4P860aN4IC76IJw3qjmekQxR89v
k6NPuJhXmdFvmvgjyVNNRBV7+PCM8J10FytB9mtZUeMf1kRZPfA3F6Cdn4toSVY/c8yZEM8mZFAZ
bt+/AYJuQey/JsozrJv1+WGyc+mASTb2xHXFP3KXmtIo0F4IfC79noftUp1d9TolZhIMnV4+fYmp
UXLbDNicjRNQ9/akZk7/OebYqqW70kmnWDcVRT82omsSYTTZ+pzfZn0IARBvozKqSc0njsuO5VKN
kLSdepL18lGkBV2J4nhz2C2A9dtqwwO52b91HGkvVUvWx57eFobL+MeQ/aaK40KdN7WPSsnXSJ24
Yzp0wQYXi/0WOJASLeVSJPln208p8f9V/YYJk31j8yj4zonprEej5CRmY1PYSHj8jr7qQ0X6ZaxS
mvbEgR5zHxVexxdzcsmxJCDxfRMFRnz18H3R7I+mZo6ZQohcUU1IMJKezYTQ842m5sYdxQfCC7I0
mhRiK/q2pCDvuiiH+yccYW8EKInATZt0SKZpZwcIUK2+GlDy9OB6tbSKw6NNpsb/6xHvbUPdrwuC
mpYrXdAtTN1rM80ivvASL6gf30nLekxg+YBTvQhM+5CWc0puJbdjuYwMymZ/WpFQ3XxiqXzkSSRW
vVjg5XiiRQD1C4a/ZG7FFyWnVliL81GCwU5dK7TlM/DcSyePH6KUM9T9aQN/ndUdfe8l7g37reS1
JEPBvdqUeOeN7ZsPbj4gBGRGRlOMRc2pbSIgulawAq6i9Ah3uL/ZYFDSR7qQ6BtlqcA7Xp8yQgJS
xE7wMrBFV0iihmyNlWTxmH7R7MhkWRSwMpAPSOu3nfTC6NESYMvRyEViyoHJExZuOMvm2qdvXckl
EcsKgjQQ+GapoM7LCkeV1pUSZX5V1b7qWsRd1XGhyvrhLYomTxdQ8jz2kb6BxufgVfeKgiLqLgm4
DF4tiM0Fco3kC99caPvDileBsi43C8FPERX/kXMKt3Of4bhdOxtilYXU78Pz9+LAQ+hjOGBdhw9h
i54RLM4rPCNw4dSQhVYcv+Ot4b3ohk/oRo+CWPZFCk76mXbQBSmi4w6Q7lKFoDmis2RKjZ0RhF+Y
jJ7y7H/0CuIxndCR74tu2MQyZvEKOrLHIcPMGRTU0AYhR8XW5CoLClb/6QFoTMoLpScqJprdPPPq
0e/U7V/Lu1/+3rtqIETiGLmBqK4lLTWy1yR+fob21GPZMCtij+d2EpE3tr8dmkFwZzcsZoVBmxV8
B6vzZBvHN0ZB+MiKRIS7xswbIdPm9VQIehsWUoWYdvv8Ms3aVEemKMazzFQrDjJJpv+OGX5Mnz+P
kS9H4p3YbLpnrCIwHDVhE3c7TmK5BnAZ17BLwAT5dmqRpd5g7q7IGcnnGwe63hvjPXcYm+ML9dDS
3ESdRdin+KgK2DmTp2bwtcbxjC/TsGw64gH4UyrZcATJxJcEBLwYNKwBeVyfGPE6kRf3FXAFBBam
d0PsViHQ9EwC0L9+twpgoA9V1PbrmhYr6wsXUT6GYYCqadXcXNR1x569kxM1BcyeZPJG3rOspt8Z
7OHK6TdMY+KeRWGaXcT/YtbQaZ46t0yiXG+V+e21ggWU7bJR7lU07djeFRYH4QFF/NBnwRmORu9G
WpfAsR/8HT1mK/fxHnu9iUOkm5niM2NSpamnXVf8n1upTwxUYAj7mqW0gWgyqC0vhSphWLmlNLDN
/qh4obdQbHoin+UvPEa+31UyWJy66OWkREuEiTgdEmZK82fn9teO5l2x8IMt9H/B9yqaST9u6t8b
+zFgAJHfbEW9x3JPqFlk/it3BZAfvlna2L0kczP9U9QPwrfZPvEYr8tzbVRD3zA6aeU5ARNEMlIr
ZmPZpf+zfkqFmmQErPUUPujNGDC+3c6BvBM00ECPJYZ3+wn29Jwr8Lkj65j4nSTNG0+3unGwtW5z
lKeSXJ2soTga2Kle8Lknl8eMS9TpHmI/1IrihkNQfa4RC6k/TJJFx1cwDmcsLgsVHYITpqqLEzad
x8wigJhpkC83Nf6iFQ/serFjZ4WWQBgN+BM075AX+NsTcXL7ysfKRRzZomdXaYnNkLY2Dxz33yfn
yG+Hn6hXRJxdOLn6VCzs28yR17Cr8Wg7eWuqe5/cF/Ebt1eKHqLYVZtRLOb2ApabGkEfQZE+YJo9
7K4/9kiQnXGMS2pF2FzPHsa4tbgCoH9jkdAgndqx+1zoMBwA1o1r2OQj0Ly/RGj6c/xr+hVlC3sF
aA91zoEGRTN4ktDqbGQ3vki5HwQY072aLo4AzEsYhrrN82f81DJ2fZlrdkBfG6ji06ZejF0DcFZN
3S4bRYN1Erifd27EnrQlgtOReWjTZPNProk/PpBA5Syvqpi9zYAPoJIw7kJ8hiIKXDaPWtVENQsW
+z2X2zR1BeeejR7yisqWsGDoZbHVx9mSGCz/bHSTU+2lu1crcfFJ/Az2FbXggnlJbAbd/UD10i+k
3c+2XtKZo7JlEM54tseDoaS2ENjbGiEy0GOj65a3x4rnmOBBHwX8ezEGFJg9FYmWEu8WB/H4JVGU
bWNZswv2QH8/Ww94e4jwaq0Qfjo4j5kdlBr2BxxyeiJcGz97ZKYu5xKCEA7nnb0oXB4fDbcLySGT
nyTwyMs3axD63ba9thzjNNYACkV+LiH0/ntNSBmxDX78aAQxU6kUz17xm6qeG3Wpr4o3/ItK70pZ
ZHP76pE0nejnRpRgDBuH5zDSiEguQlSNbEd2QXEp9Fpc1HJBHO7O6Lrwfq8VMJEgnK9jdNiJX4wp
VR/ZpmVRnyGTXRgq6Y3YS9Gd5HptLb6hnAfxYJk6c5m4TiRiRz45xz2IITkJqLYqkuxg1NR2+tIs
kxzHXlNowXNmocfTqGXT1vwcA+fjdhd7/x6zu8tTI4sdevxPB1rKu4lSZNb840yjRE9uy+qxjpSw
IM3v9jHUwZ/hjkQfuZkXHtYJz2ARMINGqMFx/Uu3Mtp6o88IOLrjj2G2tPD60toNE2LecBJ/QQ2j
Nf3x3YjDufiud7CIwBl4j+PP/UALXaGiIvHNi2I1/6QhFKmD3wpIqRoKOwmOxjjJRKmjCDmtxInf
4y6yJFH9WHa74DOfIcQcCZKgXtN+i/6EGO06JLg6JZWOj7lUCvCJyjGB9ZA6pOs1HJdIovU5UoZQ
1ROQse1rrshqNqJquVUiCA1AVpr5d+BFSmh1xK1QSQQiMy/vxRs5cWO9UamQ+ClTRlQ0mlRk5GGR
70vLo52xoPzktge2TEenfeAohKb+0sdnK7znmIYvsmLhbgvi7TtAbp/rCFI2r1sIFVoo7zfXnR7u
bD82PIDOz2fJ5MAbgsPvqcUiuSSfOhL5vZ4xVRz1GRRR3rIb/qe5BWw6ioUmsRlz7cvu3do9s4kn
Mjvoro2qfaR6ZGcHb/VcgBMQ+xBLt5jL4FmdrmqoBhvA/rAup5g6a3GLaWcBMMblTRPuFFKULtsN
XUlSm+ClfeXiHVpb0TV+J2bgLkEMLXIGhf+4VOAh88UaeIidxiD7b3Oojp1iBtnl7VUjaHwezZzx
ETQr5BywMHJCmTtdDf+xC7JiW7qJ/MvAD4BIqk8Vm796S4GcJLlp4wq47Hv/nbP+1drXEFQB2d+p
7EdPmBDSvu1NZUZde5RkZx5iJn3p68+Fj6dRncn7GY9tDULPtojifvb7TNfSlXIbPHzWDqQpLCaI
Hdqah9sVVSS9NK0A7KS7wp8KEHCXiiCbiDxOzL+LouHQQ2SajIobGY5Gx1wepkE+YybkWUFoVkYn
DjPWTv9Ud0YkCsY1myYONd9bjLeTe0/zg+ru/o9bee7zfhCDZofCvCdvzCmA9Aavh+e7XvIYf3bt
n93gpzh3Ynnotf5Vomp3JHRq71sNSZYJ4Q1iq7Y80j6kWYgWWt8xpIpTTRRLioMsuzCMnJLQ2rem
Jh5CDHRtMiprCnPmMJSCr6fSWC6G+a7klt0OLpDAdaDXWe2Ax52ZIxkG8Zw/BwzOlmkSO7JHhrvM
AAGYRfe7n6EgjpmC2Tty1FUWad1Ot5LDfgP8HIoTLiIc/H6IIvOMC7vt/MdAQG+dGKbLk+w81GJ1
Ol8ojPyyBVNw5Pw8L8zocZ/A81hXtmAcZ1D36wCxnxZDbSXeXtuZOB277dtNBtXbCHaUSrzpbp8f
0CguBoXvR9V4v0IKBPNnQzuehJPCGAZSiYRJ/CU938MiJl2TS2aG5G9ZqFpUFnBef0dnyaWfg21T
ELjTkVzal5vAfT9Tw/YB3QniGUQOgOib0TAtfRuVHgfKtu8yo2kfNwtCZtSj444GRxNgU7XYL8bK
t0qZ4pslLHQw6vmCa4aHnjWYmesjiKce6Le56KSFxtfQIAJAlHP5Tlm7SKCBnKCwJZZKoHmi6jPX
2JSqr0MP2J8uDGc4j5csGOWPn4uYcK0cKg5pA3GmdZX4pgEGAEo0FUHAgL1h4TRC53CMLYQcFiCs
YRgUsQvV4H5AQcAqI7J/Pxe0cNO8i4i+Wrr/iwK/5/39wDC47aoOcJJyPYMJEaJFJl+SgIgq6Rvv
Jp3qTPUoKHdS9MwaxGpKlmgK0VNksUBOSJyZcHr5Rbpa0yL6njCYn6hOCAgjVSKN/HACUBlTDAY2
8EczlDwovbCnrFiRUJqXago8h5UNKhRVaFbVoAo7g8CotGAsWa2SPutYKHRAy1zFOJAtA+38a7i2
BmD1Fnb/qOrh/741eL2TJGheU4tj/CxuDbaR0+QUnFjO+yFp+0fMAbimkIuulUTrp1mP/IBgvSuk
dvaHqfrDugp0FARdTJ91u98ws36qNrDw2Pc2Bm5FFNUETLWke3L6ButewObyA50pPXUK7RjWW8rq
nYQ6o1YWsbjQiNlx/4jzIiJgxcKDVHwdHRmPCZay9lW+N/tOHZth2h3I3dAjMzFeUbWW9oEm2Lev
NHGQNRTX3+kiX7uT2I+U+G2AEI/fSNQenGKWKTSdInnXWOUaxmbFAlK5E0ig7G/AnD62+l+xSxGr
ect6L9t8QUvNpAfjXFsqMOh5v43swijUE0JcFMuwd/STZ+h8uwhGy6z7OkWhMt9c8Q1SZNWbgebx
tZd9e6Rvq0y5s8MSoA0wkpcFTxI83l0QazD44X+fVbLjPJt9prDQNrrOblsyDU6yHN6IVwPFmIrR
jxwoWYDAPI1PfRc83YaETGO7XQCdvDQ9JMOmOo58DAc2EHuheUqX9uYBOb8wavN0Wy+zO3GxHKDV
dXBFVda1AZWYVEHcP22kJzOXigT9s4BtE8GjTaGM4iir6tmE5fO9mi9NYFMIftYVeJdIQ+0SRdsk
RQ0I/qAR5KWOIQ/dhh0MmgC3AfxRz2JCqfakgk+7dQ+f6//MjWEvUxuaTZWh+YmFU9LDysWUEPJI
BHuXLmUzQ2UO4UEfK/1NSqVD70Fy4aC+FtR1iNbk7BVloK6lphEGPPD0+xLMGCp0gBiJxTqWKOpg
+o86M5w1Lhx+vHGkJQW/Cu6QV3VEp/Vp6Ml5Kg4xHXO6DABcN75dvXgZEUFh4qQYNXUdbvJcP7Vq
Ypey11TbXN88vSefWPbqp8BeDBeU+iU6Nb5SoXErRtMEHeKGzTKKn0je/cj83//ugf6sV/jf4jyv
QG3yOyMgWu/mII31RkoaS0fbPOoD7kcCAAHxW6tY3BvS7oBXGdEh0s+V+PRXZ0QfO+tNwYZ3417C
guVeQ2ZIu4Rfe1QXVmzQ8JeVSlBHvwYJb5sDAF7/w6g1FwOkS1jO36v1VBMxFoPsXyvvWqGsBhx5
Op135bqudD75a4h/Ad88BCdthnU+6jYVbqxuV5M/HsjWODOoeWaq6V8mtTGsreBB/n309mHZT4vb
8dykQz1eUnzSG3v3PQ+hr/HWy5v6vP5V6JBshsGD9GtkDM1rMHGkGL7KIko20hKd2Fd8vscSxs5c
GN25CerAe1ZZ6PW7gHZUAFMhn+r4DVGFGabDMQODDvOPZTn75gAiEa5IJbOAe4J/n7KG5zeUbvON
ingWLgcmQtnS9FDBZ7jbeJa77wuVVmjmOa0ksK6qyAYtfNezG6TH3OI55GxbmxgjiWHKAnp0cej8
93rkrk3s9txMoeOak5ksndyb+RJH8zxZOC+itV5y72S1sdaNYfMX1sKT4n3+KQPiNLeuQx1rfxoA
263ISfsROLb7ykR8yzx+sX8eRG0Tx5xdDWeF/hU0jZvb6Ia2YRu0EzhEVrGSbh/trx3Ap6FKn8Fg
RtV9ziGa7UyzOQN6P1gpur8bn9/kpLX0u0UzYLt/enkRofFvGIzZ1VzdAyQRid5gglm/xdwsmHlX
wPZ5Drd8ykGGGCL3a3E10tgPtMfj9gw5zPiPHsXUecRgBIUqlb6f9tMFdazn3Lr8x+a/me2J5m2V
KMb0qFHAGtpMgNCFPGDEALHrL9IJdn17V+KDAJuTYyXxA9EMVzYKFniSgN1gQLnMD2EW7P3uTA9c
yu5rpAzV/9Bg2VP7MT3b82EBP4R5X5kobSTTeoQhY/hni3vfZkJV5hGwkWgJxw4vl7BkXHvcJkgC
vSe99+VkDmMru04+tVWpR0R6UEmcU2CsQA8NfEN6STNSix2isdiSa2IZgrTMse+EPKK+IfDs4IZT
Zo2htLvFtvzpTWH/8ePamFuIstq13fCg5Oy73qGZszJaaYndH69dBd0qNdZrzs/h1zEf8jF5r14u
ybbeAECpTgYKMYfEk5+TSTA6L5r/fThkxBChE3j16jjDc9wvUmjX0kctb2rn1oUDYbtLcJaECocu
UR/0+hNw9B1zkCsPOQNcxrW00+zfXD9fnIVnIGTyuxt8BkAqHjOKXZX6IbG9GJvw8GXRF1fxD6es
SxwcNJJCPCYJC4Vjl40zaulelgsHqYJ7K1RA4/X6nzkHGbv9bx2+i18dk9qiFX8HPF4u3HkqNigv
HnHX9k4S+HrKYWoylIJldOPCEBMdalnVNP+Zh8CB0gUrlcghN73/eSxgvE1CrvB9NYAJ8C1qWOOF
UFvdkJhjAY8oFeIPm9yevvGR9hRYfQpZ6pBgw/j3pHpRoHAybNC3NLZPuvHt8A7JzxkTWOYK+XTG
oaRtKmQ00IiVut82aerXWODxFBwxbNfhuLzA/BO3j2gQXoCS8LHtvDfiXqGe9NOiL+pRDBXwKPaG
KGfWpLMCmYRVJkuZhKuNpf17Uoyn1Hr4Mj1LW7SB+UQNJCcb0OCm4iWLCS4HJ8SD9trFlXnSshWd
xP95EHMtUXdFuG2PWIKyy31P/gZEf9Dg6u7Kp5YmU2qScuR13kN+qTK4Kz7zDpV76YKAwROw248r
qu5hqGC0swizjwszkbf8qw5W5/rfwVAwSQoZVexPqzsTnAHC7/4gC2OOXlw6wojUcPweu2VqML04
N41bmVZVtTiAU3Vg9wzERca6dP+WmzOZB0kyiUOCARJfWJ8nfVLERhkCEUBJLlaz/QBlkWeEIHTq
t7GicR+ymTWS2I1rui55eyl7RBPg7Kv5hYERstGv2YfMx+wzsaVxGMwFaz+WKETqEiM2IhYiqVV4
IYDDOABlRYmvjx7FPTR5Z7O0cBFgn+N+FL/UMkgiqpI2e9en+J97anDPrL45faH9yOMwkZlx4j17
iQ1v5yIB1QBpBU5a97vkdOoRrvmRqCRj0h8DNTNBPQG1Z2J06n1teB9tPYlqZd5SFUH+i43T3EhD
IGc5AxMYUKldCpd4aRTa+g0bmQAwPu5qZGY/upK4w1WKG0nctHAlmN/8ZciacA/3CDe7tnj05ra6
lOIK9Eq8HEUVdU6gHkNBfNaV7H8LDzX6x4UuFt7IWt+/ymlkvIHUIPVUIkVNhijdkphP9KzaWCO2
jO9jR6skIGmqD+6FDiKsN/S4i59wBnPF05Bi7UEEp1ZxlU6211R4tO3ftz1PQWgcyMlTQnwRohcu
ViK3j6eK9gvLzquPFitwRAFcWIOC+goRT+TdxdO2sR6vEs5P4w5yQHDD6c+bHckHNPmtJCij8xKm
51g4rjcYF8LC97/VUee/CByveK4A4iBkicZwLxKVnKNommiiVg9vSVk5YPEb1h32F75wz0rxZdMK
oDHQ9GK797NeGpkQiVpc5o0f/K0bzNRBeGNzWZMgBkRDS6OuSTDGiOM3fKyAXPWktDqQiKMDOE2a
+s47Y85ekZugxEbqnHK88ZoCyfCXghg1QuE9b5atIzdwihhSpx+BNlLqPdp/N3GgPTBMHJDzRo1D
BmdcHa2FvHEZ0Q0mF1VnBa7Ru5L6UBxVaX5K8Z2CIECL68nBXsQ3Sj/9oiDGtyOj39RSKaEAjKDh
LpEWd3nx4EHAmv+xNfYj1oZ6XHJ046jhCOSEWjItbm1kvgiGmVgNObtRDtZV6vQzdSclKWrr5x10
D5Zv/ur0wCaKLvpNRRNpANnFm4v074lqnUjIE/xUoKjH4ryj7zqaFumr9oOldYeI5fTO19lpTTyc
AF/MpayCmzPe69i+febaQGOJVTZE3QNG/V1MFv09jbj9mcxp8pJMYwG09Uv4p1AKCEVEvBi3n/40
ly3Rmk4uch5mYd/F3gtoBh6+vwDn5vO985Q2cumxgpFdFqyGqZc+rgxhgZ3sjJDgwm+h4ghbT24Z
RgGDBYFsH3UANMByjM+tx0WCaf4AOkzhRZNBJSfdSgJCW0dBjKa3rPRP/YNrup/8T6r1lePO8mbP
Afe6BNciISfK+HU2GU4mqTI46rkHYqnoul/mjZSfnvNtGvhTNhvSJ+QP9XNq+8/kmMfYx/thkyUx
OROt5y5IV00gCQBluvzPcwmXF65vvG9wQp8to9H87dgmIOJmy+gflkrMUsly+O86HZpC1ToXY+wU
H0w2B/wSJ2eOz1sXF2Odyc6/6TrdiSZv1mLyiXdmm6LSg1Oq2v3+dWDkSlHxqPxbngkfy8Nn6msF
fgG9Uo1v1Y8C8w0ztYnYPeIMnqHANWcphAwDRAISdVic7agIHuXC54KSl1fjt7sqgiD0CdEtm5dx
SR6oxneRB37g+pU4F/MfECo+G/719Mdwph2y9ZUDrKVd2EdEy/3vXyox16Nl6YzXHHUq6Dn/lOvd
gtS4C1LtLmdfskE7IsHMs0zUvJhlmUKOOTCjUXxl3HdL5zXXEtal0gpWBKPefWwXS3l2TfkVGRFr
0XvoEHpqXdUt/TxqCqtl9S0HdqyZcjbRFdF1N3oWtRiL1OWuSlVGkscwsqDLAoOIWbewfs6NsHBg
k9xxRqeoFh4XCueGC91AsxQ2KE6zADePM++xWfcgZcowIJU9zqoCVAVAHXynTOf/sAtHX3XrRs9h
GcInOsbZPShbubeuPrAwjFmtfOp/aa4hxJ/x7tnJ60A9DtFqFnRiDtJ3vTxCTmbmueMsQnN381Jn
J2Uv0cG6N0VcBvoe3LL/gm05RzBMkBcb5s8WmhDvCIrhO5V7nJtNedawES7eMEDkXDEZ4t/BOCTC
+zEMiWvth+u2ziugZyVy6V9ktLdMG1ktSVX1usvbc6KJlzDBdnPIsMnnNgfkxRz/QOFqagUduGbg
T4xMcV7Zp0rGGXsAowe4jGyQqhK3C0iR3Uf+Bwq8D3M5X/wZC/P6D5yyb4W/EJFpnSyn9EJ66ZSD
OyC1RssBLUDHAU49l7YR2Y17OOYnM3BRqoKMF6GoYEy/Za7SzAFdAFzTcpOc6B+1Qahep0qGt2UB
n2PjUBVHWuZJAssRZZ0CSY5yvBnOE+bD7MfLuML4BPv7QfTPGcDcPfJuE8+w4og3ZJ8K6B4IU0WC
Xv1CBcrY9sMmbuBuA1jYD8UDn9BP9mlCTVPfyAvoVcn80rRMs+IqbcQ1RJfGUaqkb9dmALAEorti
g4KDMrmeywhqAoZ3QLPN6muqkO6fkSiGp0OlguxVVSm628BLmpQC6svYuk6C4oWtd5ZuJCP6rF6p
l3i5z7kspsQ6C6JOzhntVlOLwI4cQ4Ck4IMbcsF5jw3lck9XlJFXBqLFSt01kHSg78q8lvIB2QRZ
1IGMcLgPvM6KqiZxrC7RYycfuq0wEASoaXbGs5mqyJMfc7NZ1lYW6sIfqANBgY9YCONtN+XY6BYY
ZIIrzc6LD/agUiUN1ajy7kY+jEGBev3NLLNEY81iuIksjAFk93TPA/+TY5FqB0DL/THTP9ILU92q
wi6s5l/g/2+kAdVsFbOLLadIHEfMZFlHvdsmvkcBQvHNWVk9T2qK7+hlZ4SaBCkgw33g2zRY7D+a
NCVwePru4c9YVBWOXLlaeu5X+RuQjNvLDtIUbUMNhkSCAFYSe1N5mV2Orv/7t0ceg/9HQ7oyl1IY
N0miWRqRm2NoSSFIZOvRdS7sBC9j/RnFWf0zIf4pB21sy5JCF8r9TIWn9bTWHX1x1fZEF+ISCM+m
arZHaoW2dkWuFewkd50zU6DJ/gHiJ/W6Ao4kX6G5g8q/06SWnYHZ6HWsWplHD8pPmY95SyWVLqQn
EY0sG4I5E+miImklhEjmKJkt2QKB0cgNGCn65D8xXJkM8scZkF3GS/BjgPI5/P/eZw3V4iZuF5m6
O/D5l79c7ARcNcjnhyjG1FjFJg6WvQa3Sn7qmyq5r8lqXMZwKtnQZwQMBQadWN3ayiMLJG8s04uA
saHvZ/3pBkeQ5gxixxCUDWevjfuw4J4l3LcPBhjmPQ50ujstcQglu3qMHOHi2SoZp9ZLybe85vZC
ayZvrsPvJIKqicFXqbwj4b+oKmy3jXu54ZyaG6/usERaorZ4Om54h8z5LKhizqk4OQ3vSj9GtXyN
SsC27oxvHKjEYz8gdkcuKeFLmsyK5zkax/RYiYNoUgvAjmP/QJaxGw8whP/UcWAH5wuV4/VL1WeH
PrT6CdZnVqggk11ekbk96LnBNCVv3JEj86866r+BlBT6x+h10Ql5bN93b0SEN5fx0sHlPu+SGqrO
o5JL+17R0MsqLklPNY0XGdpognyqEZdcNm7hiZP1aUyIp9XAtC5rUySwGnXADCku/NeV+rpch+VD
Dz7Tf/DDjVOUzP5mwKZQCHeyLwJw90rs0GwfP6ojjyK8k+s64k73QlVLPjrNYfZj73x8z2wnTMWG
85duZVyc4UcPoMhBw/jmSvcOr2VRa4REwcjmxP93vn7Ayy0ItIxpHDOZT7uY+Pw+8C7Oc3C2Zzj5
Hp7no9frBgOIbec5tVmHJq4XJgLqhTQ3aNQH6/4q0XhHnSyRngj/Ws1s3GwaavVcIN1xP/GLe0XC
nH3+QQnsS42O/NfO2v5w6W2RLt8p2IQRuxM8VDttefsGAnOtaEm2a8GjEOs0FvHsxm2eJwyKSNrg
yxNvIhHymIHQiB3O/13dBtCzxappiHSI70q8pJkiHsCseIOSZuxNq+pU3aDsPvi3Eoz2U6FL2/XI
CffnmfLhDmvxg/1RTi3inWQFT2Z5tbc5Wad2RWgHVoK+D3ZGTsFOpSkcaaYYvoIcol5X2bfb7vPG
VbRD86rXS7KwJrngscipiQkmeTqe4UYmm9I/R36nD4jd9NZw9ImG9TdJ9O4lltlERXCfUQaQJYuc
K6rRr3jZLvvCSbkKV2q40dxfnquIkEiZOCbfnHfeYhJTAN7YhtB5ASgWf463D+sN6PVdsAjMiQnR
zwc1fLkVLrsWlIFi7nK07h19xvb8OB2HnACqJEpHvM42G9aKk9pZH8Tv7ZC1abjFM64OlZTs3elS
+QDFLqf9KuObvvKyOXNchscN5fWL81oeVjHuu1Zp/FdE1N7sUPBVhIWZtqz+aPAtR+YlHxhRP593
gWCt99mtoVgXUf0goG510Hogz9K/HnwkG8x80iyb8PiRCc2kuwDUok1oFUjt8f1U982V6zN2syFO
XIfXh+Yk0B8maWBBW6Gd0xqvkIWktE7V5Fs9VRoF84FUDKsuqUgTmKPLcA8/qFq+kkPF2k1Yz852
XzLsGUygnNzERb03x/+Adgaoeby1NoX+E/9Z8UzOazuOVYx6ugE8xbgbtMzVpC/ep6liAElmpqDL
GPaBmeMTzUgA+GC3euF/W2uONNf8sa6YHy4JwpzY8gxA+gLLhzmZgxnObxdVp6irISaDT7XsIROo
zsPiDci1gtJEnXnAEPpl/cfoFiO7dOd7RqH7gtu5agKV0VD3PdDIHgodkSvOpPSAbAgeEADqtPZI
AJdcdEEmBYeaQsYhGrhec8fw5rdXJKIKkOYk9Nd5Zu8tiD92tc8VLDXnmpCXkceujnvdgcq/VDbZ
44wsZQEMnVEBq0ryWTbuOrJEYx8PohguNyzhZbrMgdsPPQ8W0+O8/VWD1Mkb89jAcH5XtycU1JzZ
k9Cnn8MtyxQx7vA5bz7XlXUzTPfQM/Rv5QtOglHTDC0Zwn4zDdbc1LsIVaTRCd3iYnAa3Nu6smQD
2CKhRHMNcRWWgbgF44PbBokUwrFY87G33VjR7Q7hZTKt9zu4h6huBOZI6PmuZmpgihAnhPwcwr06
lKnzb8DdWKHAzyn9Ol+ujS8f22ylY5la/ck8Pjsu5wfZo1IFZntj/k+XESAv8d1PDmGDS1b1cKdA
AaWNOKx9xXZ1CRRZq9v1UoffqMGbhbgdOSBzxGAXYwFOdSiWbmKmZ1bCIrKqK7qL7+HHY+ZSA3Zc
fMN+dV1UW30WCufIPh8gzhmQxTFJ8LG3Q0GSczILPZIavN2Q+DlNY14IkKD+DB8Ea8hUYnGaf4mw
l6mdJp1nzSPICZ0NDjgSfBHrDbc0EZ9x7/un1Dx/JTauZmihGqHq6O/bGUT82pfjsIvaLF3DpOk+
nX5a5cX2uhIJn/7bMwLTg3EP5moud4j7k11cyV42AT2wiMz8KmOmTCNp5kJeoL3xB0uPrtjhSXXq
QMrQtblp1gPsThL95+9jYdo21ZnBpXAe488BCc+ZjMClTQ9AZNotZQaRZGPrpgzyrDHXIx9oIRGh
jYKzccGi71UB3nYahxkLEOejf0WWsNiadki+pCT4tngneTYqy4Jga/YS4GPx3w9Cnhu3gWDGLUUT
6tSpJkf5V9tM42RVCiQHl7GvXmc+65ecO7hCdNKyuCoBVEcBuiL4gghhdvTGwR5Q3ljVuO+GiFAP
TFmbXx/Ejyk1IdS9EDwGOWmw6PSBBN9mapPEcGnLUG5wh1FPBP8dpV56Aj100poPy+KkhITnk/T9
CKef2BITiOG9YHMjOjD0qYdhaWbJvqt9OU1pah6ahMRYpzArtaNC8S+Pg/F7q5Y5OKDvFPSfRUYq
p1a4XlvSS2buKOhitASPqBigtKmZxYHDrSNpel2leJdN1ADWYs24S1Ogcm8c+RsV0AHyy+rprPYy
9IgU4zh9+nSnQKdj012Wolzb+SNNbvHIgm+ycptHCEo1aPTSS/aIp7ZrxfH6GxRBvSudyy1qMyGB
R7Y1JGvlzFb+dP/jJ4427FwxXIEnWv/m2ccZ96kyCZ1bYqPX8fJPSewhb8IGOPeIJx3ACBije6DM
t+L8+erE2FEgRZoIEQxHI+TLDVkF211cKv4f1L1ea1YY9KV0jgEXXJkthWqjBAurXUVTwG1/la1B
yeJ+J9FGm7MuVMph6okM67TGv+KqWrAJ2AZXfpe51BUcwlo1o4hBsGCjoe7SMfN8wEo7XAR37U8I
HoMJox2voz+uE65nvN53fHXbSpqdyt/e5AsOLpgb3eY92lNCL9oxZTMF0hECKD8dVVFM00HRIRxY
zdlxzhRTwODlUVhbRE6XozJJ0aC/i7PpZEFotuscjVq0f0eKel/ocJEg6lpgt6L6SnYCh8X+5Qwo
9aHK4QN7ttTQczyW+MrZCZqUpRee230jdu9YwwOvIMpFADk0Mj0KDw1KwJu+7SepyIDb0A4eeGFo
4DWfaqRcAgJ93jWXwm1xxdOj8TUOLq9KL/bPLC3M1iXnWHlsI3lh6/XKrX29T7abZdlCNBCeQ7hc
D2vvVsutOvTKLssF+Llvt1oHVLsp6kGjbn/vLOc4CvNdJQH8K0sj8VRWrqgSL5/7fyYSLA/7D3mK
CgbWUhZvVAm22NhUEPSTzdcQVk503eUCbBRrKIbtmJNmwuNSEab4CAre1uzNXqdrfRLZAygq+/XT
Wla/NrTSFpmJwDDcD+Y+aSLC8pFFyGL0IvKbYfmRjAR5c/TofDI2LPuZWrVcvxt6bSfzw4LFzwRI
ycz0O3KllRE4LQkU73aoaqaef/ckm4Fy3ejjsoSPirjhBFtWMQ5O134igyTofiZze5MMFU9grYAD
wKt0k5A9J3YEcmbF1D3ugtnuHGYlv0x2J4ZeCoTyLdrGHeD0fmIvUbjZLoYwEuEpIjDeZHBZ2bDd
TzuOy6NtpO2QWvbFsSp7ae2iT/cowuqQFNM+t78ReI72MxjdJ5VsVp0gXGQEqlylL8CQ8/tMS9pr
biAe8orX6S5JEr7sgb12cPGZFg0eiCHCVg3CKTB9s8EicEsD32mpag7L6wzuoc/P15AV5NmYp1be
ejpJEIrXkZXHtBpLbDee4xeNEbcWPMfB3DDwwzej5oUNbp4/mrtLx5UAG2Jf2m01diWj3OOrwgeb
/3O9cURAHbQwqJSqo60MfuwdAzSrBsrQxYiJt8+nBo5xZ7yBmSdd/dLy9HqVxy4OMNA+8g35KXbi
oANmzbUoSfrC96+sInsc0mmK1/PwstAk4xMqpK7OhGvwCGR4eOyw3xhfWwxkzCw3Q3B7lA3+M6LF
ncXkGthP4rpBCRj9hLP7qyCQdjtQVZpA17OdoF7zgDtM6D8vOlW9BObV4qRtPeNBl9KLL/TYBNh9
SxrPxTmV+kxaLw2vlZQUZr6vulmuNAZVx2D+25cgN8NLHUyd24BX7O4dmtDC1DAoipD4XMvI8YYO
rHctyX9TeAj6qN4eAi+ieuFzBt9ji0s6NsaCfNwnFtU39ofA9npAgoN91ItRPK5ediLXmkC/Jrc9
HnbHs+DJIkVfwzznwVHXjIIlnxnCIUPhhh6mmfOv60+lXL999VCyXJpXEtn5FWAwjdGuf72KmYH3
yIIEeJ/tWmSZlJHq5I3yJIQ26kbftjfyZ3HE77OWQX8/nXQNlTQomBuk7GfyXk+k7c898/bPN6mm
L7kIVF20+2NQxcL680EcE18EIpYJ1QGFKyTpNQ/vPccucZF/+V7dUyzM1wgkciPMwInFNaYuDeGl
SzKkw99DGkcMOkM0vdi6iGSjfZB0g2q6Na8fuNcuGgXveU8X+Q1iITD2wjOeCjSlVrEMW/jZ+l44
aA9D91fgDcMaZVNkKLvSXwHlfC8MhWMV/semSI62dMlupJJEt0Mt/rn8dvPnAh520lqWhgD56mNm
20oCx6Dq+W+OhKZmcOa1bIEkyxkln2+E+Q5gzf5XIQoICp7xXrMdaHEvZGHODHBd6Nsici3egUXM
e/a7y77yRsNfzjTD88QlQNgnsHdV0i+0V5la+fZJ+zxdFoWZPL2TpKmO5+kIghLVHX5GnrQrWZlh
jHCkUzFoaiavblCE5cflCTUrpI0ZR9xRYRB/8idDx3+eQ5sq6OxMNXLvA62VU3Fx9Agqp/IXEIcv
2l9Fq5DEvqc68NHsBP8ECK1vNSC+YIm9ZTgtJYNryn0LshPL3OEu4yT55pHMAqRPFW/b54i40Bp0
bDsh1EQMlqucLfHHjzm4b7mtpDnxoFAi6E/dh0iXVrDCVDFT5TnK5N10LUDeXtZWtniHAnMYdxEZ
zu/eNPCZVchx6bKNU/rXAQs9XMWkK+cN5WfOLG+4DhHILsSKpKVGeeB63kAMsPRTcJeDkKqF4f98
fiI7s0xTNZ0jNufis8TnpjwiocY7kwe90yg2cAhbm1W+jNVWLYj3TEc6GGPQgX544R5V2LfNWesJ
p7hpv3eEa75RHKMBs7BGaK8CNJJ57vD9j+d7ogI9SQonAQWPjTXPRcd0pJE8AhppTWv4yqE2bebF
1Skhh3vtShewdEoPvR85lVMS/F1rUiChePN1JV5Ii3yDa9eZdE9/TEvO/FE69/2BdV2r06TwO+m5
ExGUnhxp20WkI7MADL/wPJ1jdjPfMEH4lEYp6kNNWaSiPKkdNG2rH+1Kr4b/OKMLudmd6DPvSaKY
NRQsdVgPQi+JGCVN0p7HLuegHyZrZRYAAEoY2Fn/eBkbuS6FF1MTef27MXtJ0jWCeDPtL49fTBk8
ROYMScTP4PlU7TOG0DYo8hkV8LnhW/ZhpMkw7D0cgn3CYeTcj/YzBiVUMlwpYrGbrJDuueBobDNG
AOYJs2M6kEoIRdj375qX4N8zO1rL1RR+ERcvUi77rVHHVddSAXNPgIbyfReEE0qnaQe0OkAiIlFS
563PKNOKsU0/qb82WbNK91OZbALN2ipa5i5Hj2bgsmfnAGsM0EZpfKYq/ooIRz18wl1UKXFOMnOa
QvBCSfhxxsJQMBlgwAnTPNJziEMqlfoPfb3vTv7T3oOrIsi5xoZV0+Cjl4C+jxJS1dbHciImnO50
NviRmlt6/MdUTcrV39wPi0B3t0HFJ6Rm22ejuCl0rheym0oNoamelh4HkV8RuIFI9CVZfEKXJpPU
sswzqx1haYkCrSCy/QP3T8BDYbnVQj1G4JLh50uJBAhDOVxmRSsVuRXOa9jahgF1PmnTNT8NG9VE
Gw2BjWZBUWwDc3BSt+dIl2hAxelGuKCPxMx1CUmcoMVY4XTJb3hlWQJkIgczdQzHyCSJdHYfyfsu
bjGUsmhXjfNF4T9dXsPaU85dwc7nIvQ9anfpbQZGj2L40ZbCY9YLXVd7SuTuw0JerMAauaZLP6W+
/hTRjQMLPFHOHL6GfsU1Kn/ug7rXfBicz4YG794baVbUD1FjCyvKOdRogiEhijYgHpUlgCBqOKjY
qL+gofZ8y4zyS6K9FpBDgQ1CiYHlahjAe9E/fGkfIX4wEIgPoupxs8O/TOtPfbJwFan3RrGQypUd
0YLf2nsaz5LeM3Jhd/il74RpOuGM/5dv5kB85W+b7ZNDZvX8p+JpczI+r2pf8MNUJ7MxVhQggWKF
iZw1iSDZZb1v0spstM45hMDJu/1DLzLuw+guklL1zZVjAi/WJ2dGF+HMnhVAJ0DPywVCFdZRMzRw
C3qOMkJs2/GMEoahVidKNku8NhMX2lbO9Jmkkthn9Ort945d8W9cnMumUi0Prt+dsEp8lqF0L3j9
Jg+rHCHtXkh9NIEH4yv92zL9AnqfFi0QC424P7gIdekbCyz0EVwqV8KjvlOb49SPteusWYT4m0l1
7mPpNcxk2oySWszvKRVv1d67YmCyNQZH0R8RwBd08LbFfqioxKNbWvIgbBn2MIBpigDuvnsn0NSb
rs5BtOH9tl36pOl/WOtu0rcXk5pazonlA7sbAenntFUrE8p3KxjFddp13iraTK2oDoIUE0RKdDZ2
mXmipB2QysgnZWZK5FcTPcITK7qTMr+Wo0yvGbBQT7y0nGVlv3L0oa8wWMba+bykMxEPHVaRjKt8
kb3yY/9nDa6T2PGx0wmNHB3gL/VjOY1JYsBCx9cs8JX/Ve5cbey+5MaceATUlUEQgwDD2WvE5Ubq
vFDYAHS6qaXdwtWjBgsdCRY3fzPcSlXk8tIjaiaszykw3VQoNsPBU2HsnIC2ufMDHqHMflsRc0Wr
f9PZFlxmD6o3YVes7v4pStrh9DG4i8wtevr2PnCmmJoxObF74499HKiBQEMD/9fAaKOoT5eJflco
Yb03S2RIJlFMvaPb8TxYWdqq1qQGR5N+QS0EgFsG2z8uDo29zy7IJrVqF0SLIMjdPzAdAGAr0RKD
uSCyCLoybCPTbiN/0tgVLul5A0qp4q3hKAGfa4W4UBvHr3U/83P+HYblZeFrLKVAQyq1CPOvS6tE
TpNsyQTgxyuEpOOazDMwl/fsiZlMKLTFuWlvompKt5gfRWzSlnuF1e6ceYQinPuHDmu6LdvxNXjf
z1y//ClZR4hOR68pR7hcKsT18wNejjBGIiyuKfLu62XDYxOmvz4FlhcxfG06RM0cMtJ8xKSSQQWi
BXIwv1AD6eIff/L/A54lQcB1Q6+vfBqsNkAA5Jl0jFrjbRdcc9ZcjvFY0LMung6SN/aFyG3Kb957
aBt5gM6Z4YLn0CNYdOX9Tebjk2SGfawYcbv8vFUBAveuSr8k1TR1WyuYgRMxX6ddDzoghnt7u1Mq
BwLvgxvtRgma7/MBJKSpk5U+aN4CNjcDC4lL14PKvwIF97PdSiLmSGDfD+a3URwYUNYHpvfnSFOW
+KwPlFv4bcsufJPkpqkEHidsFFe+DY+xPzfltq6WM9c2l5oYHAu/KsOIRnvK8Y2MZeo13WG93ZA2
0Kp8gh/JpVeSwASv4Qjf/kOpMGMC+U5lFncMx1qQhsU476RtS8us/ru5ZTfL1MhUkgywcwj0dwMv
TzBRhDBbKaXCNK0M520CzumoKg2re1DuRENKr0HZa2+/rdiv6HIlTUEPcHrvRwf0EW/3DymgF8aW
l9SGewTdcWMo6OqWdw5c6o5GJDCn3XtQGBcP2jX81z8rvmqJQJmarufPMO2j5pOnrzV1BviYerJU
CCm4kOXQCc9pKPtiMpJk/f6uY+rSURDC0dNkTMCu9w2qyHY+DY09Xf61IT2U1q6hc+ImU8NOhidz
quTHB2KbWFBLomcf2uVvsYehOMBasnMWR+UpQkM3bHIHq0HH4XrtsAeH31azBuwitcy3RGOkxZhw
7YgrM8hdMo+02mpxEl0rNsYv4y1y58ldKaQknZch3Vd2jw/AG1d1vle9Nfh4JRO9mQXfpa2l18pC
8Jkkz8pOzR/nKkVIghNoB42JcQXZZrSdDEyXIJB4yWI2fbjUC7HkyqqwzpACejOkBDg4EKg4nEZ2
7J3Y+GA/VkxIt2tVy3d1A0JXtRYxP6mjIarHB2kKHnkvo0oDaDbvb0KFwEakNulUBGfwxJ+5uXSR
UC6zxcI/PsyGEBaQIJ+zj7srxi6Avl2K+wnuiiRE/G9VyuROSoBkPvhZg2T0WHJc1o5u870w2+gM
x7fUDSP8AczCpnaf+VpXJ80O5JYF3gox8f1yVCUInV1hH67jdPlDHTlfrg/zthg3TukAIIaTsUmc
Sba+dK0/w7nOt7UtT7tco9vgF5ZFVkZrmMtwI1gGgF9mgTAMhspHOE67Z0n+1keiDN1QIDD+txsW
C7jISIghKgt4N24VxmbLZBl6Dg+9bixQ8JCV/NfgCt/XhMhElviVpfwI5C0jWL3t/yN+/1ugprwk
qMc4x7Va+tOvMsDS88ziydtRqNvmHJJloJryc9pQJX391fef1aOvTs80SzRNMLQI8ea3QJsF61JZ
MDJ+XfLKjzFOAAYNEXDAJeGm/X48SuyBXwao0OV5mkMo5yZTOSFqOTw1SA0EzxwP9/QVMQ67agkI
UNYLEL5D6wqgGaWqwjh+pYt3ax8MG9R/M3RDwsZFSXq7YNAeEOhpd+P3+Mv40W9KPd78LrjIbKQb
jxrm0A9yWhochTAyaJBS75Oc4Ipm6fmlZNqmVUwtGVN6LRVk5vkn3V9TMpsF20pgXN5/jmfD4GlY
bZTacU3QtGMS6ANxE6v1knCI1nXHzywyKa1rXpkLXtm85lsD0U8ZYK2H/6pJgstJhZofNqIvQF2V
TNJaFmFtf0vm+FTFWgj7XhEKpah4JMRPd+/wHwDiSfHQThSNbNk86a3Fg/w/vhvdTd9XlhJCIcTW
WwEPxQnXLoW8ssw+lc2b7cb7Lfw80SNt1E/YFHlP5zBaCGIekxwqqwrmlGsyk5vhlu6uDPzFab0X
ALQRjHVi9a6EpVQa2gfheT/F3KVlrhtD8q5BGqD1rHMDlEnSeujQaAYjLp6xlzjjeYk5OpTVPbXa
StwTnP+2gL+Sh9FDHzs7m8ZCqFJqQIyZ02k3EWSnbVRYLGQgI6CZjMDAIC+Fz9+bspYyR5VQPgJf
siZJfTRHPT5ym56cb6zqRngsfNshN3w0njG2JCN+kAO/5RDI4KxFuXzbxKyKbFWQCVbF7bAX4Q3l
tBOKw+tq8YNQG6tlxlrY0om2fUR0Qv5iOLVZnQb327qLQUyiTdU3qCFxAXp+T/4bS06zduQCV9k9
kBIQwcZoKpjQXKzBRlV3LUQ1+NPS7W9pUxOZkuS2rPMO1HCInl00R1EHtMAVhK8mhPo965tv6ArU
l3njt044DMo97bk+sh5A3qkmOW3xS1pAR/ydBxO1+6zzHS77ga/t4eK3lq8f/TkvCzTpaKqF1qle
Q7AM+q4smcl2mfVod4VQsaSksqN72FrybOVTmy3cGAJERmnHIR0id+2QKpayXXPMyZp+kUMIf0Bl
ZcZywryxS04ejP5illI7GpmeHtsRWA/ODqJSMNDd3d9ZAmcQ/NftWJSLeL+7oH5GZLrAGtuJZMFS
kJmfxSD5vBXUqrjyCZbD3YEoooY4QdHWEg95Wn9oVoGTyRsV3aK8QOlyYrQveuPba7d1PhNQxUbv
hXEzp4TX1wL3Qm/i5JEUu4uRsyEqiXizztQXbteKk5mixrdnpAOruGoC2a9Jm8eHyDDQ77QDbQ6O
1yufKKn9orHT9XvtblD1rsuedvP2UXBM8+B69RZhVlzd5q+OPyPKrbhPwHd59U46A0rZXRbyUuiy
Ha0YfEZxzGh5ZsA4stIaCJORcBy0nfDmbGcT8EJh8wl1XCbLsDa0Uuau4NDQRwLQUeFoGti8PYQD
4HpuMyI2sUK8wYUCWBZYl+qEdzIy6RttlRwq/w6eV+LUZVAOTud3G25QQs4uGcSKLl3XAXgoB8+L
wn3fhC0Pgj2eZD+dO/XdR9O5NUSn9VMVnTnqsnK8RKlM13FpBBB6+rwXPa3+QagPGqwb1v9oQAQC
3FfHvwRDSxCklJPQBMnPyKoeGC6WGuM9LmRTIlBIpOx7Eu9+1lZuKki9xgqQWPCw0nJ/qgvse2UC
1KHT1tb0Vy9sDZtrBdEM85SGC5bQ1sUUjS6B8spd6OSMWuIwP5GjSwbLYj3k2KGBrFT/EFQzmuq1
TocxhErARXZ+4KUFXZ4HufyaNAzoM9zdW+Sln45jG14BRAAmPGeVOkMr1CQtgQAIF631Z017KESl
s2l5gMFBSlH3W0UWL6Ev7K4jzUTYK8ZOFdgh3Es8Ah88HMKdpOeKKQILU2yqfQa5SK453n8V9/Qp
rKmI4yTh2s5R+TVMroJCNW2ArZgIdeyRr+0W5WpZzRnDJnyGrig1QicudvHPKHEMIXb7P+zTOdy3
sJsRWzDeHKhTfmDZUhx4EoeYPQhdBOo/ZUUTxNFWrRNwpvQh9t9FRHOr5HMBBX2MuVEm8jmxS1Kh
Rf2l8jmS/lLldRDvJE49zzs1sbbz/sIknYtpIRacbJPvco90xv2TNURIaKpS8NCTdCQgvuXVyfdE
0U7+dM42mUeT6JnZ58he5ED31gwyfD3wBPci0WSP1RXgBSkDuZZKMn2RBeWEDfTOAeZbwOQarazk
pN8bjlkpORWV+Apq4xEa2cJD12+6T4TNxCKd1xR5inesmEFbUY9ZGXyhvT7DegjZxuTlrhpQPNvW
Bk2m9gQfEq5+nTgAC1DiA+hQBp/yrBcgi2D/8yb9ZrxSjoWg/N+ZlHKxqMgPPknS6si8vWmN7Gwk
Sx0EH4plhwIl5fmnTStOJLbx4XLlJ0SmYPOtk/CPDUbvrt1MhBmsWr55nrRIA13uXYXpiroLYpq2
4JENPKYVGEFo7vpTsOpaZ+BraWMLZ+gY//O/ucLsv9jCZm/NOTxcP28nz+ELHtWZT1lZkgMbFmHv
mDYTp8h+enVDQhiPcaG8b7py0+2ReQwEqcF8XLtZfcXMswKnbkj3gKG2sFG8qVpcHYBMeUVjGNam
vXcXhe3q1Y2d+hJoHNErUwxkT8z6eOaUIkcWoOoPGXymZ/vOmcki8sewk3OX2gAe7wtGrNh22vny
tb+MeKaokpgW+fj1FVYN7twivcLtJ8uIrsam+/rGSOYmYegAiUiHQTCLLh1j0JQb1UPzckLiUZtW
agd5paguLFDR9a0r73xI44lF3nBN6DMQMH57YUlg/XjEF9+LgGbnND69XPpCF1U/xRJkwCvnYGhF
8zK5OssJx7TJdaIVjK7VevA9Sskm2QEO/uDIYKePs9BEZgeQLXENjcrZjyxonUNpHXOrlJz7SQDJ
obRf6wOFBNuo0cQNCz1LKPMw8ysBixFLim9qzf7Su4WFlbCE04Sn7Yn1MFeq6XPmgBMwbZWfqUwS
kO226WepCbzizdxH1mXVWGPs2ie8eYQgJzxJdbpm4X99g74Taf4PeMdkwoieznwYHI1Oo+erYpdh
Sb53UasOBuA7kjEO2aAE+RmCxqHK6JZ5bdafwoTMDnGH2IPV24mhxjQL5/Zz8KPc4umMVmlnInpw
rOrFMsnfKDIkY5Ipp0fcsbQlSUiBRnXTOle1Bssa6FHTvjHLRaMxWoW6LhXVdU1PEf+qgcSm2XA0
VZ9EUC2B0nphknT8rBBYlnC65CBwfnhalX49XnOJbk3fCNLzdr1nMPxPb3tabWNMFtOL0zs9efQi
jQroeYTC0rXEeGKojArh7zafqp5jDZw3CMJ6aNAvtinBD4vFeu/QPQ9ruRqHzjNoQDLY0pKY3pVO
8BdbvCDrB1obJa2sqdXr20L6npRZ+THngGLDy+PzBtrXwhd6iUlQ8JT0tfNeSJx0LPSzJR0nuLRs
jJxrhX+tk8euRLq9donl92xBTkPy1LgTWgb84+lXpleQxvMNtFe6iPjc7HI+2ejHRloxDVEvjE7z
dlzUI3Zxn0g8rRzeAh/rBJ7Dw1AtUQIvyVwDqPC+Q6Ex1LtDIX/XmKEYst+ulK/5llZpNJ+y1SHX
8BrEcRzA8IUrOI9kpjIv6dEAK2o94p51pvst/uE/lqt/YGGMAulBPvpDjvwURPNtaPJw9xPXK9NJ
VSyGxkK2qQY8NvS3eRS1csL57/R38hlphl1Ak77lTtSjbMl7iG14RRVvbkq7SloyAzMyn8kyueQ7
2eMp6qBjcQzafM+zPRuEreWSp5SuIOx/ew5OsrUN291j/avIvduIVnaZADW4CNa1uEYKeMVGGPnI
N95R+VYwtwpHG+LMGSHias5C1hT8Wz48pTFP8eSpr8FpImDM9f7PhLTy7gA4bjNUIZzkvUFwVA1W
G3iMcAlc9pkMnEt0j1yWc3UZo4n0OyHmopXQktSENanv1n3hYBR4jywTCpdtHYxMDn196u6IgLhC
YPUXU5SWDb5hh6PRqyWe+tnsc6TpfnFB5DUeYg26/drn0+1XHRlMIIP4Wk5Ru3HBWtfbwebLTtJj
vlQpFPUGDAXsN7iclbhs3vdJq7y4wssjBhLQsyczjOvfBtZs3REx6MI5P25oYLf62o0nVVD/d0DH
A5rXUvOwSpbn1JmNU4FQ925MyHrbxRJBfWFx/FBwN6LQeW7O5yWC36mzR8FRNymlNcsFxBVzEWUg
+3Jn0jutmx0PE9u0cGUBzKmiD5VgudqrcZ0XUiFT4VIN4DnqebODf8TPws12t95exH6AaxOw/SHj
ubtp4t0lV/T/wnJA1gUhXiI/E2QM3jYDGLkZoE74GKVgZeInPfoNCBNYTcE4rnE5Nh+CKtqT+bDw
w0fMDC5JhXt33QcguoCJ9KB6N409JTOlv0qcE/tu4rn8VYRvBtWcQ0+I1KYaGg9ZI/4TGGBgw7uG
vhV71iyJsl0EqXmg7Kek7o60oMoolvWY6ZUjx9SrMFFUc8R8F4xpN6jAOlGt1kRuT7iMMJ9/+RJX
WKdrZY2gmOrN1xb9hhz3iCwOc51cNmP8u80pm/t5K0Q8neAfny9IPTaeCRVCisVEYaRfTpBRgU0v
RDO7xwllPL69NgU1GFnPDUDrWfVjeXFjtAaDjSa3Gk8Dotab1GPHcEuEWJMb8mBKARjL22PAVmbb
wSaCe4yvPkdICerRPkiovJ9gcH0BJp7bNKPGaYaUuAHcQo6lQdlzcbS1p1yBFy4PjfZEodYr2rvV
6ZsVP5JFi7v6V3wvt028gp51otYI4s6Wx6xy9KyCEd67F7iyQwh0WjcbZEu/qHe8IlFwMAkcCAmE
8azjtEX+Xcv/uf1lYXMUaYt/VjjzosiwzmFQJGOe9a8UVytdls72RsR03phcWyONGhGadItOdyVe
OyuQfi6plCmBbjs2bWUAquioLILmgV5ABPZ64ovCuWxHS7yYnvyGE4GKHgIypzZyufnsZbdx3DMR
yV9xIeLzu0IXHZpv6/MSerPbYtQ2TtvgfXjr3o0HSmyyp+W8txei7CXWY4CiakKeF2WXBa31GLzW
JNs9ucE6QiyWvhQhEvDXxHEsuh/k+5F45coo9XvjDGUpTPbKHqDoYROC30t2Cp4SBcxE/SL2K9h3
jKp9Zw4PcP1S+5x9V1lL/vFNHFmRj3PbiSSEfzP2UEIKr284j5y/dEr3nsVNCiLIVBcCiKCwGhmI
JhjH2FhrY4s5keWlBknIpi6rC4ssCez2txhS4DaTDy0Zf8TZEZ3e0XzfJ3fYKTPD6HTQgRJvm9hz
99km0xw9U9uavr751YTiXluPvNzQJGn82xKUDK92RGD1rm28A49Y8JYMykQxWtzsekr36Yi9yUHy
DjKVonLdgpNfpiTf/nfTI2Z064wMqAS8JweWwg+vXKFVCQyBNiAbRlgBHAOhgQUgZHy02j23jZOM
zqnU5c1rW1I44tWaM+3aNWgq4SJ6HBYJ6WsB1N3onlZSsUL0AIW4wY6LHWwDLssc3R1jEyQR4sFg
ShZARyAUBaLVBvcoHGuKOxiy03xV3gaPo2JqUjVAV7kFKP7uVpNRZ8ax6bbeAoC9EtkivS9hmBIj
nUtOobrypqzKrlbsAmQjFjlcMRM9Oy3dZ/6/1q4GLDb1C7cFMGhA2SOXi1rdnZtw04fZSRQwh1Xd
/jnAY9fr2tE7hQe3Q6YNQg3kndg6yfx4SQj8zUqR7GVzMTIB6cYF3r9xAUuZtN2hsyedfuFZG0Po
lkFjf0Zy9/0VvvYmtYzVcndEWKv0tdm9ErU8WbltUm/HrS9crTXaWkExSvjZ8Wxhac6JXirU28aD
pYXPiz43EbyDO3wKybsToWHbgZ19PfgtCXK1Us3ucso1IpZbgDjbCyxWsrHZQ2zlwPpAiLpH3Zyv
c5tGHLK6pyPvDR1p7AV3dAz+FZgJ2TTCaU5ZgZMNWERPjw8ECzbzYdfhaJckVk+4lDOWQGfauY3D
kjgzkD52idULsFzIbwEWhpRcpOWsHdqIvQqySAfbqD1ODxtinhUKM7tkjoD8tbO6H9/jaPqZKKHm
szdRC4I7GSsIwLU5tQD2aVZOkxUyA+CyNw2BDflWyn/WDBPrWIwp32uMIKeCTOkr20I6KERQJpyP
szeKWllTbG2IQQ/PLYE+g3TPX2Z9JQ306bOrhxzfLTN/PpQn2HNmt5mO2Fm4/azPCiiCq0ud2gFw
95hmp5+X3yUdWNsDhOX6zFGJe5csQ6wmIIkUwFJ33m+SBJ+JxlvcTtCEfc2lpJ6Pgc1yRG2yDbO8
OXH8bGgncf4UHNrr8cfQAyfAeJKBcE7ilb03s3TKUonKOqdLLu7984mAs7ZBAvIGSwgEqzsEF/XK
/KOS0+uwCK0W9IP7jOWP16boRMeua7yhq9h9X1ZuZbclEA9nia1BqDE+rAscEPc0jU07H2qewjig
imomSh3uZ44SBL/Ork525J1MGNIQ1/Aj00T18aUTqTKOSOXjcp9X0G4W1CI+ZtKAhEW82yweuGuF
QhGTVmdGLnfZvCWmzpeW6MqvjLDMdEBW5vfFvsZAlvEQCQey/mMS05XiiyurqskkzQgovs1DbWty
eSNF2YtqRn1/5uoXtdZy6OlUJeMaDK/cxZM2BuIyAh/THkYeoOE0Rm0FYFIspe/bxw4Omi+Sws89
pAmJTHxUsLUQtdzATUaRufEALry/qiZzOjvCMBGLAAhfKWNAIYnsATSdt7ePGSUTSP+Y1i8gyAcu
k5TH0qT4P0UJJTh47yHtI/UmriLPwua18TmLSXPI+AIL64G0i6So9XfEEV0vKAU9/U3PsQDLdOQX
glLqTKb+V3RuC6lZ7z774C9x4K1o3F7WPlrErOG0ZeiZVy4xd+YIq2GTi3n36+fQOSxXPbhrZYVI
dhDyre53W0sshdG6D4F2TaGUIbTgf5qUIBfUzp8jtYmzEGZiyMl1SEXwbIemYFUPzArY/Fw4EPU5
b4bxmNA3Kcaz6ojccdC/IzT1qlK2cLzdquPEsfnVTzYP7Wgrjb7JmOSmQ3ZLFc4YEpmVDy1vnD97
P0eEtlWbT+BJEmmPmckC+uX+GRs0aU0Rjp20FSkTBPbZAAxFsPBCApc68if7BJlpQ9weXJ/aPNkF
ixzRvsgJbCZuNDL52bKNQ9i0S6iYsrzZlWFSdCInuDa+v78vEIkx2baibknSPvfhDFURR7XY6jDo
galpPc22GMeJuki3Khb3bokjjKQeHedDwq5OjjabwbU35W0W/D2TT23C9mmfV7M/FN0iXxbrNGXu
V9xB8Us5vrC/2A2P5S2U/MzcBwum7ykYjoOW9m2CN198lyAm/bemz/xstN2g6ylg0sX7UnOgST9p
AsBRWHHKV5uAGrc2mOTXZvgMXZGKHSz6RdpPrN5uek616z7IWRzrid6Mx6gNnYUdH/cZuCxQg3se
gl/YbJWVvfNPnbmTFRGWAbXW+PVBmLgP5W1Vkh2DVieoxOkEzjeSxKjAeTeqnHRFE1dVarKU7YAG
wxrl/xZU252dUSfEtSQcCW/M2F3QHuLBrOLr6M/tg2zsFazPjAGFuc5wUHII8Aq589eU5bW7/WGr
1V8A3XVpJMm4HNscrLwjgGqJCvkch/UuWgedIDzZ7ttKkbTDduGp0C04LNIBjfAM74RQM4Mpxc/h
1zKsxdB1Glg0rDN/+dmuylUWpaqH1tSCHs+5n+fX7lQ+Iq8jJaMi6jL5lrLiBI09/Jpp+lZWoA83
dgc+fg053v/ujqISkQ671XsxDzBP5Iak29OOZV/AgeoYEKH1Y7cNHKQiDomt5MyQo5Z3v1gsKQos
2TZQS1HEexf2izPVjHpkUCru2stKGWts7W4cmpgl2JwyBURMxAR3QPGfU1AAjLK1YuDGW6jcFnNX
4AyjI83vCV3OH8cmWvG9IZE0549saRO/08tvMl8MFNsddyYHU3QamQaH36fag0Nz1FJAx8l2/B8t
LcqSo7rfO8vFZmv3Mnvhq5othN75DXZvfF7+KQsXNnWxbcLbEK3NnEbjjaaNIq28sYI59NleAnau
PDeO160BXgFwFPZwhiO1DIxD92QGpPPccuXLDSLeyDpF2j04xhrtWmy33FET1ziN9pPr2AdF9gGE
sz+4VTlJWVwWqoWWmsggHAbvETQ93q0/ntmXxd6h3u6sAGgMwJhE5LD59xc/mpifmDF8If7diHq/
b238kjGdIfU43dyLIU1mCYMjVIjYpqfPqQh5dPHmg6az8vl3uDBYwDuWnya/YpWlHSmQuhf08q/3
YAB1uT36YAkRTRrzOBV9ydUBUDDPSsXbt4pRI0OrhwgvbuXpoASnaYBDFi6Ozkq7GKKPQw5yhZca
k8eqJXRmVJkzJYYw0hxijZeDeRJ7Nq2Coe5OiJtY5ac/KCLAz1ecfN1MNmiIelYUesNWVwDKQfRu
ndtMfvcAJtN8ugm5zRJKeFYE8TyxaMIfhAetusaMThajYcTZ3U6grWr5y/A23nUdaEONGPg+EScF
niOa5fY4m8TzjkDgD2erzgYzlRrUTfHMsyHkTRB3BGEP0P7LOjuqe2+hndzZY8a9gcyKonpckkJt
jrsChEPQ1cfzYqc6G/REJBrooWTwPPU+6QaNPWg6tkSbNGOMYohNTFZ6L/ygW0vMja6x2Jc4k51l
yXCyd57NBQQ05ztWthUMRyXmmmRQLkqhBc2udnxk0HMIPbWT3S6jPgi91k0EtVCenhhQF3rz4dcH
dO6Tq8MFphhrJXRoxMHWIQGFep3B0+nei/ttCVO1jqmXHOeTnTXWh5ZpxNrnyM/tBRfQfk6l8M6K
trODm1/vmUtIOEXJKE98AZ443YaTtJ8qenElJmr6vZNTpfegvIXrRyTNmWk2IyD+nOuuhF7blVbl
oqz93j4jyIDuCnPffaniuyjZeX00cih4Ubg/I/RwXIXXQUu0o6j1MjoboIkXwysIsHP1BwmvH20Z
N+pbQf5jb4UvlDFwMJaDyfvO9k427/TGwi1QVDM2zHCsSZDa9NRdVeMtRFz7dDMeYGN1kVWgxqdb
+xjpGxRnsTBXaHvqdNcNdMI+REQmlC4tpnwhrhdfz0SxqL/WgeLEKg4AAkyqgq5sgVo1zFdmgE7B
Xfs1LKqPriJp7cOSPmB8yyqGmz+ddilkiTWdzRifqnwBAjx+a0TIdWLPLGKUArSXHLS2yKPguWIe
akLvq3n/Onav3njj0FO+ofxdRy2F0tQGheDithFp0keog6Lm35XZTHSe60OuQv3KNHWDSBDNZfej
ji/LfHFbElKEwDDnCqEe2MhImturvkTQLvJX22kuoRjJkujA8n67rCT34u553B+BKrtV1RUNZLNZ
xTpH9lN8HwQZOzah0g62JqOTJxq5ShXSvdvSSNg/z0+fk1hnTAr5psmM9l7s+GXBEyhLPEyMBlwB
u+Sk2nGpTZ+ahxOq157+iSqVCDayfaYRuBbx+D0SS85ryEV1JlFF2XrBykonydV677Jh+85hQT6M
k1eM+IgaNZQ/NM9mPPNVo0ssXQQ2TlRJ67RLNxdFcUlsA/C/HftCrp2pm86B306p8rG20Rx/Nytz
jE0c//hTCpQI+AjppAf0QC+lbNbTLQkb1ELxKfKss7XX4WCdI/1M9HMGddgqusg8O0461V6VZhET
k11qq4bkt+50PKNjfQ5kRz49C8v19wnr7f5YbTsPfqoknVPWUazjdvHBEIJqPqXsJ1D0cElpIVWN
VQtyjUX/JPIuVkPXy52M8htwux8deeeSe/e8vUslQ1ZV6UcvygFB+z2vrpHrIBscBxqylsj1woQo
Eg+lVbAIW/DvMNwRcvs8X0omJCTaSY0LqtLR66k9KCd8GhKbojJsZKqHAgRtV+LZgLJf2Aizltxz
e41gbNWNHsp30Is4ztnLUPssEbqt0TJVRtRKNi3ft3mmEe8fhBcV3EbCnJ+HdV4kMg4lQtt2/1A0
Do8/pSxjGrKp4EQ9Kwzmmsg0xl6rgmnk7YLURxZ/9khr6A8fZ4gsmwqhU4YorLAceny9BPAtWaOr
qEZSVgZB0AuYKMNmLxF4VqCrltRSeaXMimEp8zyzwqzDfZWJO+FdCIP1+RXZecCSqRvvQAm8Vaen
scy2lEajskHkNLCXCYUaLMJ/+sbx4AoYES8nqNOb4778cSL4K0jX1WIgS/VvkQCpLcvNuokyDwCT
S1sFuG5RuiUfPLXVo0J3haJ+kxDo8GMtl7NgBE9BeGJp3v/5da37HtBT6iD3MBL5leFNmjzOBRxr
dnT1lN02Ljw/5/VVSn6hkfuKyYLXKotp0batnyK6IIuaj5lLigM3YmqwQZW+S2A0uZ+tatjMrrjs
xbzMffRbPImXjk3HJz2iBCVlY3DrUrmya39R/GTN0/+rnvP2v3j54zO5F2bNPs//nqek1CPAJzDR
9JG13IdNlTsOSqe23C+27/MvlC5g57W/11G8ZyfoQ6XwdfBO/mCX2yVHDGIZqQYWySYTeV/C9F0x
ml/+vVr2YM5flMK0Wwb8YSnSNR/+Zj0CDqNDsdEErGrb8Wj99MLp75Iupz38YHmzcwI7OTmHJ5Og
z6uNS/azt3l4x0SqYGAE8Hul5S4T6889zwD7OhJ5RJB3a9IobdFLIeceGy4COErPoLIFbIzj2q29
/Pfw8bnqU3yf8l7BDDqkmPKwUJcc8n51WHK5Hx7gkmAM8GA6vCesWnZQjDHt+B/xSfzDOmlk7V8o
0d9SeBXQpHejY7HTZGNurqHsGL+TOU/zRRfe9jv6QQY1EkH015FaM1ZYijf6bQllxvQ/btBtbfMe
wTs0mjYwBXPTi0CucjeD8mQ9GoFrXwsZiCwkmuG3aJj3Uke5EIN8oKMgpTC/wXUQFrZA2Po0+Xh6
6MestMmkrD3Z4UMgYe8czOurPVh0nS+SSH6Mta1TXQwfhQVBu8w59QN7xluqiYDuTzY3SSBBYocA
+PVJr0GWqM0igrJUzpJHE31WnQ0wawwSg9x5voMwpJKtL12P23Wt5Qs32yvKhg6PnXGFSfDHaq58
Oc/sWi0t/NtghQI4xBr+wwZvJWL6Dp5brw9OhmAsCp97OzKpaOCjOAcOkUPPG9Cnhxbn6HrpOCrv
sCeXfyAXdSSVnTPwBjtw1C3NT8rQk3NtseRyekTPKVxklXQK5fwK76QULTwtKXTijpPxJmQd8tup
1g1ZBnhY16++oE5scuaCLLC6PMbFwDuO2KyGPV3Wa+svhs1irFXWFvC/IxRsco2Fh+rM5Bk0gjE0
2S/hN4ZBobhL7hshNcSiNRxRrwM/wTNJMEO0PUV7IcfEQwkbyBScCrs8pjGLw0aUJwKuDM1Pp2yy
edshE4Uimf3BGyynabtsjYAFbRlN1mPJiwRX6QrReIxAJ55dmkCTVrc9UrggnzhjwzX7ak3xksHP
n7OcDzXvadFwdGG1OzOEJpKjWpsSSSAHVwn1Rmftsb5r1yyPnrlTtg4tdN1WccaC1S796usYeN5E
g2gLjIMFdYO97juvpSnlpJCVtjmTshdfI363ny65WR1DUwqABIus+cn43r0WVMUryzp/glCPoMAI
bxqU7CgFgN8CDXtPD5Hs5nNwvs1aN+17WtKFAhCc6Bv9pW9IZ5sIj9QrPNliXEjJKztAarjVJAea
0NhuBI4CYJRWMK0ztLU2g8Lqn6478l1ybAj7bPcEbVjSRJ8T0tCX22n5TuPy/hSWPm9ar8ZGFsNY
F22RKbYiEz0elwtjp80FS1jgbv0g0je6nP8xe6Ztc1fjIJJsMv07mJ/UgsU8Rvc7MT8xeZAAbmYA
pNNfulmGUKpy94s4OVFzHYpvrj+XvsRgJkDOkQznhwgdiQokT6V1MLsmVTFkX2n5tzLHrU45/g4A
6/MMqWQfEc83XNm2Nr7JmZUIawKT+j1LrA+VL8BaTG2G9xfP3RZWWpjQi2AZ1rYm/qRg7P8nXXXM
4e/SfF/NX1uYn2IydcXJ5oV6MgDp8HL7MZnwUuWJ9hgsBoeYaiVRXQmNWm8h+us5ySq7uAFpoqwc
gLhBgkaAb9GmA72muDxJrS6FPhSO4y29y8YJvHjVFoc21YZlm70NU93yX7AS6+ogMyy6ASPrlFum
VHqvvco3a0VfFDSnN77AE1b9uxIQl+zFP9QclowqBe6ajp2wlxi7t57UXD0v/Dv5kqq+awi3+YEY
CUqspKdnOOQ3gBn6SbaYQod5+uJbY+0QMOFlhVMUqOg6GtQ3LX+C+LM6aOXSHbpuJ765JeXkPB0l
OdZtijPid8jnYaAChmK0IvybRiAgnI/CLTyq7AfiG1HBNvNlYpZsXrNG+sTCGkR1J1/m/zx3K2ef
/A27uRDWnH1KHUq96PoXyJC7qh7KjfkvSVbVjjEEqhSDRQhYentmnyXMECZSd7n4Cl3+QjiSenaT
wBUH+0WRs6aENBk8kT6V4a+6Hfrsm0EUilHNCBJrOC4fpuXnKTFFFq4uW/ztE15IqgaWrvQViExu
Vjox+GhaAU3758914JJf/pVgTd651uR7ZSUZiCvDxGXyEDQimtDXtCpbV+U+Pb4X94TiZ4/CDDhB
f08PGO/XrCDnOs2nUMMUlI1RmyC+jn44BlJVNYmmPsBdaS5AT9JyohB4h7/pUT6XjeadoeGCiueE
g0269QZMz1SWfgOeOkVLLkaZnWCnV/agC/VIrrFtgfEqudBKESbbpo0vTRQZApo8lqWh1GZaeJuG
8BScQipCTXPpHflRCJNY+NrO6XESu0j2XOAgz1cr6+EkbpCuyWcj/UVUNMO6CX2Hr+ggdyBYfI4a
AGapmbuEuJ4HfLvVlim/HB+K0VDGQCpRATs18uA/1vDXSEgn/6RNznehHenahR/ySkVc7pAihc3W
evnUNxV2aDkv4iwOiiXggIEjo5negmAp7s7NU0TdD84YbxBeXy4xBqvLq6uAnHhNLo+OhpLpMB4C
HKxAh879iyauZHQHo76ymJF6FU6aLUDi78NvpNCEwA4apD5JEGAcfhKmUAkFA9GuCYwACfZIfNYp
+wXSBdsFt3gK5sosJpfBQ1LoGhRHx6I5sVpL28fY1xLgbfJKMLGtd2F6YveEf8fmqiuYCXq6uvCP
x5m6T7FRcG8BwgRtQZ6FoUNzyqnX65K4ZrMj14FCv8SxRTwC/tllx4Mmk2JhlCInFU4wYSGxNRPy
tP47w59jkSxOI6LZaOHQPXab73uyDratPiy5QQ1vFoBGjAbfHoA+8IPeElYQZDKZK058sqAlaEf0
Te8kflfZYMjKIZY0u/KAycU9xuMvl5h9UF6hEyDASpgfE3DT1UL1YEivaSZmtCZ5wF3g1RHtwkVw
eW9RXKi3YZUDWkUmDJ7FHCSshM1NoQD6if03camWfji0S3hz8FMfh74hkGSJZPjNhIpbX/99kIkB
SfwiAwyHAK3SvyZFCzN66kQbkXCDl8mVChddnsQbr0nL6DkKlgrPaQMtCctapoP4VYBU9SM6/oYK
huwnwgWxyoRu/DIa6L0yvWtqLseaxYyvKMcV8yau8p+p2oyO3qUIXzFUBjTDTYConsqQKFvyjVjl
jHEK8NSDSP5KP91kM79kXO2Wy8j3jGlxQY6tigyTgnIx6G1YJUA8QNRe0Eh11heCU9fSWBLOAadf
k3/YAYZBDhZgCixNlcUoHzmP8QrQJkCRcY/fyjQ8HrPKslNV37EOXW229UDv7D18RZ0Yc0SsG2SL
uUucYYc0NW/vXz8k6O7/OcQT0/hsp/XqI469DjrfPnK4AZyWLDjLbtgShJQRx0+l2nzSJ/7Dg2sY
42ICzhEQPiW/sd/8fjKYHHLK8dD2Ud6GE9dzusx90LHbM85BEwC/svbLaAGCkxcWfyitX+n40hoV
64oRDUWli47mQiQEdsFJPB/FJWXlcyg6pbk4wrjj6z4pDRI2Rm1uN0llm0tMSRW48hhjjeYHjYVO
zFA2xT39gSMDOi5oNY/wZBCG/aZQUOUbjnuquxeCrwZGhoBTaaeVGs/3JFFl+ePNI6vz5BqhnPmu
8qOoTZoAGYJW02q7AvdgtJaGsp+hpdMfCzrii1U68vE52WWD1tphkBRI+tn0Cr9AmvC7sz6DpfWE
CNyx4olOJktRxIo7rFq0I+W1HpcOqgUZE2RZQWnM6xO8Iihce8MhRaYDahY3bcHY6Wc9av89dCO9
60Cy+2kIgkGN+rtQBBiX9wC6zaKDRzuaNogIKh7XPBZzdm8LEoppS7Lb6M4qvj8dXuvK7muyJKY5
KEWewKyFSEF7ouHUQnDsd8f8B5Ca2fujYQ33M9EETnDdYPFKVBuw9tripYvAKIaePsW//AdOiQQ7
KJ376SdBWh7Yn2HbSsO8dQy40YRyHtnaXkkpW2NGauo0xWLupzBNpABGlrVZQPtdk+MHg7TxAPPH
MKEIj6BkJAAcZxisH7nk4t+hV5gkOF430uhoo99zuygjZZClLKhgZujMKvyg05uHK1AYGqHI79tq
f46Sf5Y1sD8HouwdNKIePQDWKmZf6cC/MU9WAZPTR+z6fXRnTz8VTyhl5ZHJkQQLQXxz/PgxVdUN
M3SYDkarrZTAkty4cluhfzho9pbbjOdMJaIP2l3DEOs5HYDcFCRTdV8o+XMFbIjajiud7AbL8GXk
tIJ1aP82/Sq/uK1SqqgtFu7ScLJyRviZcKQWca7A7P+fcgEu58/a/cms3wnxW+rRtTfU4JOQDIA5
YgnWlh4epBctARwb40g+bHDVZgkvFc7N9/VKGoEbWOU8mwme9rINKuQnv5cw3zy6P47Ab35QP5nq
fZUxyxBl29SaWtCKELuaFu8cSrI44mT667L7GjoIk0p2HKaKqFSIUcg/ixKfEgy1PIFovvVBqDRN
OG2T1BFikmF2C7BEs+juqdANrEoN4RS9aZ5YuCng0rM0cylQhrB5rOEfGcNgz2qD5N+CHHl036sI
MBkiEDLN6xyB+IeMOUGe3X+U1Ow8WZ7kk1k/iU+qS5dfmfokaTzhZDlpT9bb6Edir+/MAuFibQJM
Mq9/AiYuHIMFfcmaptgPQxZXqdyQtnmS36zGOqx9pN6rSf/TOb2GnOGPxVS+rAUFZEXGEP8x+2Z9
Tq6RsGS9XHZ4lfuB8L/40HMhjcAfyVXreipejX/VJaiEDugEH3EYaiMzMOzEFnN37DyB/bKm1JAv
4bAwyrNQUi7yT2vJLSiWGOjRPm55opnNQz//U2z30lrxfdjwVAjXZSUfH/rGTyvTe5SK5WzDN0jO
ZNnZwUL3nSh7ny2PgGBI0igmr1REoanyoXtjqCd/PfUbBk4oRMIkisJOnamYJjQ4+Ls5FeK6e/V3
VkQEfCg0WIj0FNeSyYamkftJ0SwbESIhlL+Z9mtn2mdrPr4+wotogxTntwRawIWFeTIwTba3Ja01
LdeYUMRMKpkt2DRM4+2ajwVG2cHLPf5ZWEgAPT6A8rMOAV+iW7sv5I64RhRfGFnkYJj1Ejp1vnD0
424a4FGQyezCngItZCUQ4kZO6qI+83Q7HAiD7lj40hGXuZSkbsYAVENqWbSuC5m2rlf4gS0gWuOq
JiS2APlBzTogpNgPPsjpD2toyfQF88LE0b12Vx2sv5ohawH91vaNvAsPiQXx7jgbqor/r8GN6G4r
j24QfxRJKFpO5UpSG8wCIoB15LszoAISR+IjrqB9lE/UldTFyxwblsyVevb9rX6RKfghTz0HC7x3
Fkfj69JXoR9q6LIB7C7dvsdYFKMTc4SHTQykRT0yGOKQIc5x83Un7GnHez493RBpWo40igzTRnWY
zsSYYl9pfUe1DdXqWRgdDblPwfWsyxJKQ0h9M8sV7khIHZUoe8T5e2BYfASUg2osMeZBHtSYR8VY
U9LIxIm1+RU8TYv4PKHIB3S7qX1f+NuX3GMibTqvnY+eyPOq6sgKsa7/AbdRM10Ixrz18NMkg32f
rHoGMF4mxyPgT9bA6N6JdPyyftctchTkKE2Z9C5PdfWWq1w6+NPyNKMCYVzCeqNeuPdYUe0l6UXV
RX3PkJ6LZQwAilJ5PgJkMsCTp9K9Ygv/EgAUcNAcKuuMWaasuxNyg0smQUC9FFj0rSH1J5ZELR0Z
cP9CIhZ0+BiybNy8QjEYLne5No+plSC9WddpZcNLswBkMr2/MmpXVIkF9Fsof3QotvNgCrFmBg1G
HfbYi0jXLhnTxtZdmbweauq0d3bDX+D+GWpb0UA5lS/2X5V8V6ODCXHz8pLitCdpz8qTLeahxh97
fZ0twQNJvfYZyRP0yJRnd/Am9PX1/SvT64sKH1SuV6X8c39435AGyko+geHq4AzPhTXBPeoPRYwF
WiHEqpmP3m5DnxjZv07uuIlAQDrMFdK4bJLt77ngkBIjo1sX0ZVXp1LqBrt0sDF2S8uUnQRmcxm2
MV+F0oO3eT9oCCx/NGhIPwqzgMkhIpn+fb1ORs4h5RMMVr0fOa2u53Rv7pnB87VcnoWU+NH11wwa
oNYraY/PEm2VEcX9biUcg5jO1MOqHRoE9Vy83oYG7JkIWvLTtZxG9hY0f7EC/KzsirZdKN+qj1JP
e5pCKx5Kng/HtWalZ/3ODAOcCApPoqBiydWjLPiu2VPUaZ5aXC/Q6ZCVTvcKHr1wY9vNTFdODAx/
0xGOkkKwmuyTQ1yVkbcSNmocwiiZXvBQoAsqjuRnskrR0HDA4FmaPcn/PHq8Xkqg1W6Jlwqavyg5
ki18AvUHQtKn6TX05/jWlrYvT7C3llcqnSiOAI+JTZJQS2AEvCOoCP04zbTT75mGw0kKgZACs2uf
5H4lrE/j6yC07tG6IXbJhWzrgvQTTUBum8NtVy86uDSECz8v6EyuBYSYJCcBVLLpYJxdcvb9hH9v
iry3w9TV4C5hpSloPStTKYvUONnD5CPmvVufzHT3fl0XYGH8Y7fQXtjY7Akr2H+TPclaeYN5BSNe
9qsXiEk6xNdo25pRlUyKtXxid5OeiNI7ldxA1L3w7CswKmCOZEkmiXVBTgK97SsVofoMg3h+33JC
Zg6uT9mAV3yRYeN0f+WV93E+AQJ/1PfpughF7qvJ5aFF/3CcYslckaZyuG9WTKzDjkIahkWxpfCx
b8RKBeadsyYeBPmD2doHEZbg8xRaMcAru5lvSFiYKYHPCTKfJpzLHEwl7RzOTdIdHRQSdCCiD0Oi
P6SIPfQRW5393bo0MQkREACpvv58AqMwM8Ws7m6b797v84fmUea1itz2djRax3/Q9TI/nfI7uPgl
4p1vtlhAwlqoEjV7Q0HUbZAqHpCJu2nlhtcLBZR/LF23GqtBd5XMtPpcotX6t/AqUFQiqdYVCYx2
hnvNp9HjtX5PuVbchBaIAUMYs+dKtsVFa6lMk8UHtYxnK2K/elQ94ejHMaB4VB7TMJRrT9Cs5NLL
0zYSPzZ7YsVUnjF709Lxzu4e/ZiLjPPfvus5oT9Xy7sPeKetF87mB7uvYJ7hSnGqqqlBll/0a4r8
Prr6q//nxQqMwLmeiZeSnd9APB20Xp4PykZ9+RPFgzyY70r4W0xusq78d+nEYc0BrCUxfB1tjoEJ
okuharvYbt2sosPBSkuf9J0aqhtUpJBbLYYQsTRm1j5N4g9pVejhs9f8vziYw0tT3x5DSYlEJVYg
aVa1ppOlYs1ALTfPPzA8PjkiSMlpSliLLtulUfQHME8ecMnDq6peG2R2PnhRdJlUbrOIZxsjZECx
lD+e/Vm29/4tk3z7jR0PmOjKag6ox5Is4YcpKlxbAFTxz+XMYAFYVRH2CWpC/qkkasxvjOgfA7EO
hi5tk1Kq7DsFV+gpBgEAoAUPyA6Kdy0Xf8QPP69BYCJr2wqFKq1DZg8GsztQr/9ESMKEmfNYhLlD
f+dMjsRtmx3/OUearrpaP+vHbFLMu69/FvBAuFSqdsfwhtlh7+osXGQ3OdKo1H5NnT1+dvBP8w0E
t3vPQMChJ55Lhwlo3lug4JSlp0LuBgcfm8Rj1OPoONkQUxd/rwZtZw8lssgFu5x6tFJaYi/QlTH9
8tAVi69zvMmeUv20yN1eHb76kJ9jGa/0jiKMjvGtEjbtfe0LvIuzmqsWTMZgyh7LnZ+WL1fZ5YXg
ppCNNzQLLHVDzMk6h5mcLJbqNcpfGz6UOjpFz5TvCxhoF15nv7IJxIwXz1NikdHgNsm6im5jbYMJ
cpXQiXr4So3crXH1f1CipiYNRbOYZl91v8c12adMPRMuyZCPmxkGAtFP2l7hPgZ42H4wo5BTOrff
9koTg2q9ibmKZfg5UdS74K937lfEIX74BM00pJ3NWPxYLZZ8awRQaTcJpf3mko6b3kDGtuEZxhFH
JxmgoYej4TAQv84xfRo4uFPpNhbaCaDyR2ZeRnMWCv6m6XdfPT2H6qYVn3Rb/eq5DNHOghB2sXym
iYVFWUAYZ1wi7//BxHjv/CjjY0LJc7uCkEYqnvI5wowb/v0TwmTBViPhfqZIrhaKVgoURhotVizW
ZTsq61eihqfTunWYAyvmTYbWA9FPKVrjGCwZf1PVIs4mpxs77F37BA93LOxlpoiz6sjUkw4xLf6r
kOChedVDA5qisJtl4h01Cn4U6CdWall2qzkaKQz/pt4YLC3Zhn9CtYFl4Ngj0DUMNwReeAav/HqY
9yg8sfaQBQWyer8qNnZP1fB8+MJ5GYmGXuGvY0v0hCt3x5t9yiS2I/J0pn20toVrZKa52xvR4hh5
WgxuAVZj/GT28PnAXYmCWTfX/D+cwsTfaNGcgaevagEO2nBit0qVxtqkvC47q+trqyMGK/sb62as
UWvzS+8C/kOu5H/NTCoz5KG+B0G6XzGTa/eexDWDWMQ8trnVDMo72BXdxF+QmJG6vFVZrBDpjbie
91X1MysEcCJ094xelgi1gPjurQ1PJRZ8IYPRhsIXEz7tKnkMZTIaMqyAlnPurQWsIG7gvvT/j6lF
0hA2UhW4JcP5RberpQUKZdMmqe4jI/fznQZZzX1lvCe15VYnHtJk/Hv5xd0tQzf41/5rWAwjRyqB
Lgfdtgwptzo1bsChYJOzxrSiiNIHOS+1brNnh1YtJn9kZLL18yVbfArWG59G5YyqSAKWaKOBkrxo
jNbH5oYVDeXouVrDBr/WJoaaX+LZLdqINZ+A4Zcxkn9FNYStow40aco0VgliEqdtYDRrKT+bliPu
K+HdLQTZcUtcz2z6t8Ars1c8EQTbl2SZbsMgakUOBFM+uzI5/GnxCZ370ow/FQsbYWQQsIKiEFJf
aGbS4lzYXC6BjGkFdaVhOfPpyOJjjTFOjg7JvndCSogehMdBEoJuzH6ytn6/GnB1zrlBQNk58R8h
NTbpwOH+XBkIf/pfATTRW25B10SNNz9AOEwI/Q2VbeRAZtZiMIDVF9n+LcjY7B6HhoxQ/BA/zUe7
IQPJfEtze8K/+Tu/sKjqauCTQxaieZoE1IRHuUMPtWomY0xQCfwFykN/VhdmtI4q+enunc4tRfhX
99HC4ywffaSogHMa+uZSfFKFdmmNlWjLlylpxecHDb7RdHTnqtu4zreMinA1evevJx+f5scP/rG3
Rc2EgwCWp7zSgaHHkdPhVJUmNlrlRK22+tvfyhUGtZy5C0YCN5Gss5ZviNjbn1z7Wc8tb64me0VN
gyxlkzyAQRc00SHxULOjTDeaf/dc/iD/L703gcvr+x7jx+yf0PuziOPyXoLj6cSZNchseSpZHor6
mGAVYE7qY3sW1hII1z3NyrptglazOhHV22D6OP0bpuu/JbpfnoaZmNUhZGqybaRI6YZr3AFnaYyM
EFkBP2OzvKZvkXrZe/nm72oUeifltvdIr22MlJ74kMXGpO0oSuoNG4JEcc8mvK5OJb0SZWyrNAPI
GYxtgeVZR6glU8kKCqkJfN/6wcqaFthp4n6MwcfxEuWK3IVAjTy7xJa1gn2im+5DXkIljvj8TqhY
HkxnZX6WkzIOoeJYtNLvYwaJhVSaVMy75PAL0OUgldpK/bDfNAkletQiShRZYRMQuNTXiw2WHXsc
wcPt9N8xEPwjYyZH01jGyYvMP//w0Z9g+e9G8Cg8ryjTznRml7IDGf5x9DwUkeNEAXrSmQWxDTa/
YV6cQpiaxTEad7qzolYfA6u6SqPQXCHfGA2b1xx7kybPkQuM+cYRr4shzb2g3R3rC9DYwfzIfjlS
rvyAM8iwaRL5CQi/KmczRzdL27GHOrFn3BmhEyv0h/6wXFdlB8b86hwxxViXLEwBIJzfX9Rlml34
3UnAZp9roFBN52NZ94jXcliPaBdwKF47hkKjhrrnd8mlPuxtTSKmgI8veOdSvQe3dKzW0/RfIFL7
kp+9P6Xzhvkg/tdCiTVnW6+/dWVWhP1uT9CBamPZeRjG68kStVqLWDU6wzsDVMsC5N2VehNneoK6
ZHMlm5IjYOENMasrC9hRnpxUPTo9hbGXe+GfNl1appYotivneMVefR8SYI2j1YxgytvkSJB5wvWb
7ULXA54xVq81GcM6v5e9sjwnzavgJvLFXMY9fxrHR/N4+TqJbYh1kjiRjqUmwpEWI9I1Tal3MD+r
HgGctz7BDffanl4kL4SiQFTaeUIYmZXUSLActww6vNagUEjHwD1Z+VG5nMSXPgqpT/tmVTUBxBIH
azcHqshhUbFQOEi0U03UljswDKjklUMuLeLP6Keu/cryk30D4crmx0tSFiW1UUi0jqi5VqSt4rny
TKwNhn/rdU/c92G7vyjda++IeFqU3rKtdeCStnJ4RZxZ3nQUmJ+y4lMd/cUi1MfVZF3oZ+MnOLxB
apVWaKBDD6CDy3dU6WWBMg1CQApxAfSzfhfCS0/oxPmic05TZWMwS67YtGxEpucL431UMOw6/NN5
uohvVNxipBTLVLQL/qBywzGq/G2dsB8qf1DFkgnlNmb4DD7dkKDG98yj8CHNuS77ky/R143QcJ/c
f+peYxGPqT2Lx3WThjYOFcMXnzk2YxUc5DK5sFWEqcvV98fv1f1mEyKxrmXsw58X4l2mskf1VS76
9cw8hTb+f5+YuyCNXpwy7o6LFWVZMbIazNAyDzmogN0FRvf40YztcmXsuAzEhAuTufNPrsNIpm4g
kNuebdw27PmP06d+lZ3pSKRVAmwcGFJPf7awGBXu0oTpaO36nTsqM8drVcGrGwTlkK3Gb4cZ+Jej
52M0kvy5NarQQQghQ5dY/9ZM/d1dyUAqeFHWXZWy89T1pj1zvDEEv7MmvA9ghMMi68HgqGLAw9Zy
Ho0BuH6Xt/zJWuLN9rrbJhwwIeElYBa4OiY8BSHYMgxu84ZTl2BpLQ8hQhGVHbq6Ho8JrfrtY274
m7IUEe+osCDT1W7OboCjhJgzF7qD5hnvh7vDawbBG3MCIjc9UKSLoC0vbJCu+/1Pv5q9n/OeKlLa
RVM6G9s163lca8uP92wbOpTOvHL/uwP+r380VRLjAqnd6lqzhoT/SEacQ/frVI9enxn0lZYjhp89
9TRTRzTO7x032ItqX/GUnyNKh40WIJU4rvwlXJodDuKkOewFvpUlaxvqANY7vXMbanZG9ZJA/CXY
FggfDyuW5YMYolyBNsWr028qKuJS8GUSSrgyF1db09j5tYEQtwgC/qPj/FZXlDetBUvzgwY5ZpSq
X9K5GRGeZIvt0x9fyBtjw7C6pr5ZN4ab1p2oCKlQ4x2xRO5ewGwjXUphveUahVtjCiYXJMniFWY/
g9JqBRN+sRDRR5mkWYYk0ROI8mCggc6py4SbmgHG/PPWGgLwyurhbDAZzTwm+v/sODewr0/rPrbu
R1rfC9xVq77UJlmPkJwc6cmibd8UX0RB8Wco/hFqfvCBDZcsxxszKxxbwMiD1U0M+uBBxMIJVnsX
Ei7i5/ZNWwMeV5Dl1qyQNEvKrbddbRiN+HaTYATZlFRUi1sMggeX7/l9zp3b3Vwjwcb+fnY3WON6
Fi/FTYiJl0XntWuqseVPDtJ2ua2i+89tyjShof2LSIhqdum8nEebJoT+aY9GMLGtVhVSn/qfIdF4
Y0VEfG6wfQKHEPv5swJj7FeAf5xgIUlESI90H8bmPSEQlpTzPCd3Mc3k056YL1fYP0kIOTzqqcp8
NQv1M6Fp8aAu7Q8tGdMf6bqCHnPqinorcbsPC7g5c6zy3jIab2jEaUgcKWLRnlV+4MPKNDGL3zdp
B/WmBGJdQMIsri5w2bVRZ9w1G/sCzO62UZ8mhAWjtZRZ4zWR1FZ59ZPCf5sBb2bIWXHiqTEo74AJ
n6KsJVEaZw+PLtmLhLzH2YZ5sdSIjwuFuClCoUTsWqhZflfPSP0ZO4wysVZOlL61d8quXr+OwOZv
M506czfjRK+dPc6mtjK99FSTfU325PLOyU19X9ZX1Dbk0cPEM0YVgyBKj1DEYxDXApWd6z4Pl2d+
vjzytRsWx1tAWtw2inso6ZCVxDfDhB83d2AFHBWN9tfNUYNWvxQxdyVIQn5z/r3YTM3NZVQO4tmf
yQA5k57zjsefpiZMNA36rmb7IoP6EwCaE3XA0pjuPKgETh0xaqHsrOCeK3Lvb2KRMxNvRGJAnhFg
E+gLi/TXdHv+sbnnFrh8Bxd1QfTiaMECZmh+wDw/BPyZl39pifmGVD2rMfMuCG6EbDKhlIEk5CpJ
2IsCYeplL6eG2ZY1F6X7UfJG0d6fEsyHAV41HSmMV3IGOWGNiuFhelcJFCWsirATKA1Wi4GvNiP6
5MOnWNdP2B4jK9c62ri6Q0fsdyjHqTPcD0kYRkLq6PaqCT7I14W9Tyx8bY1GH5PZS2e5ggeffpo1
J24Lx0gfmFisSfcdBBLza9IuJRzE4+Dk1qhaXsAPhZFj7rf6IBDeZ7b5vISboFqn2JOpezfL26um
eOwNl3fOj49J58eK/GIko5LTBCr9bpyubJ/2FLVDUHrUbAFbwWGThAyknBMD7XZlqXPu9dgYFEpH
HvYuWrsWeNzMo2G3Q0ectzY2K4KbB9BDy0GT04xrTgc7L5coi8xl55fJxYhuYuJIQetovoFxKXLw
eEy9etnQcyVhuKAo5ob7yXeI8Elet6WQeKapZdtRsmQaWE/s1LcAHUzlmuyutieY3et9Y1EWkuF7
DDofOzRboCRl2fdsbPmgrctxpJ1EQNfkC6Sx46ZlQcQU6AwSAmyaft85qOhnXVJtr5H+HmEejf6S
93UOow65rTTF6Jlw2o2Abt3LNNTR2hhVJlDz/7vWiHEOqFv54aU5Pl2+h4eSR2WzN/1rP/e584De
YHmZKZkQqQh5yf0ZaWu8ZtsXVSsa97mwgEAEE5OYixM0fEfqkT4FawlZb0Z6pztCUV007bAJoeGC
YHa2DQzNSsvPRpkXOrVPD2d5zts6iVml6DpRdk3rO5Bs71M6+l8ani81e+ziFOy/Pdj+aP1ewUI8
LWuXRgX6BaJ4dMngA5tgv3UJ02F/xuq9nRbk6NkwHnmkMh1Jon6GRCoez4yAClie4TH3N2+GJWbU
cZ5rRuzLhSjOC2M7MQSNxUa8ncUM9q5LiI72HQnPDLD9C2v2TcOEjyJyOJYzaB+N0blw54T4hefH
JOwV5BdaXQyr0hWaYFJYxGPuJS/fxIjLFH1FC7sOysBgZht3cMlREzhJlJKcxEw86DenIolBtMZV
FMRcJ2eURYf1dYp1GpQBst4ELg4wAmQGm5PsIZ9pJh3pjEQeFOrfWvR9zt/8buZv77JDpUUuCyMO
VR27L9/9uWBV8ebTiNRJJftzxWTXH7AKSmBnoD0hqKiBqm5Bajd029KkipTJ5C/PFF22CxXmuTQi
76G2pZCfhu1buIA0XQx5UV0tzQpo8hwx7BBrnwcG3KNV+wO4i4jFVGTeJ2HUQzIg9/Ngc84Q76Th
lUmV4ztt+JE9VCWCHxjIM+9vCXz9YL5mDEb4MH2NSBRBTe3np39G6ar0rAvGh8CdKqUoVbinyxGC
a4p658prazvUTv8SRJwIQUBX/JnefFbppXdUVGzKfAz/HXou7Jidw/QRd6BaO+UiRA653DlRMeLE
NUpV3Cvv9QH0wFSTndHtpbFQ6hyh0Oy3IT1hjejNj3mIrdm6L7L5z5ZEAPnQauZPO/Uis2jLvN7v
+I5/5p03OSyIubZBdKPfnDcA9ccGSqAh81svGzXlpAXjY3D/9wlbNXJbvWPkI4/EIXrh0lc/nbvW
Jj17NzcKv25oQMwhS8ip2YjOwVYmt3Ft76XVzV69dmFJ6sM9Q++jvA8AUxXC5HLYTkPfyXxWPBOp
0SzbR/SCpB66ICUQR3ULgA33f3jnWRDVlqUmxkc2IglSWQGl2WJTlfxrd1LlhKdNrq/Ob5hedgpO
tsP6/lu079dYqByCjbRubXH0OQDx6NSafdUkUt27zxv9qy/4I//8YYtO6iUGf5CoI/2NfuTVFMIa
Ylz5yGR9/lJwLpvNOzSc60JyOcOMuI8QLCzkUtbgLxXfjQ10bU76jHUP2X41QgL27dEvMmgQ3RmO
6WDYcvya7+aDOyuKAMYqywRW/Kv08rEvtrKsTA2iJjIR/nOr9wj9QNU7AA7rgxUFsPS37QbeBWS1
g+pOBqB7Oqw63jQP971mMMjTBXf6zolP7BKa1ZlUKF58ZCQwSwim2OPdTfBbA9jY2r9yumS6UduS
rlAUkJ6E9atlC5kTcpT2b3BZNY/G+awkafasXB/GHV+lkSeKJpcTyZ7LinI3EFeiVPj/Dpztqss6
G5Vgcsun28W5SQDt26q3PkiWiJFUqjUerP1YcbnckcNjLc9uA2ycoGZ8aj7+Ypjci9H+Mqj+sUGU
foiA3sDf2ZJSNJ2Eqf3nbWD0eM34YYNjgMNWp9uzVRp3w+U/KxLn+/Ubpmt1B9kUh0tQ+S+CHWbZ
SePCCglHJTPmX0/93LNGzqJ9G08a4HaJ8HHJmPmBt/wDbtnfcq3anFCS3jXUs3sQVTGxYfdWcQUB
3c8LLqmh8g2igSk69LrNBl9hn3FfTld/gv3U8BMe2CVsL0mmUKtpBmmMXXMfuIRgRh/FB1vKT+x6
6cUSkGAmUDfFHtUEFpMI1l80tcUgguu+aCje54NBvJe298k3SevMgC8BxHKiJG711CeU1N0zZnKP
UH6aZ4xGNedu7nYzngFo6c6VMRAeVWulZ0dvqQk9ucyg3euUuM3UJZ90wyE5nt26Pq7X5IY5RHQy
AqUHR6PxGj19AeSVAsLdBTa2JPPMtiirdZEFbuOSTrckI6PvL3XBt+1wrlk1AwU3wfHdgjH4esf5
jygGk/cNlpwFXH8YefX/cCIaGq/5N6ExUfv9QFDloKjwu2CgDQNb3l/Wa1BAQfCYEGsSuSm6BJVg
MChQqmekS526Av2VtSLH+oZnXmre9w3aipiSqYOvVj11DQOp6n0RHo6yx/9PRu+7xmpSpWN9qShZ
FFDF0UJ/yEDx1fRHcxQujUfr1uMGi4/QMdE+bQDix3Sg1lBlbUQ/WTM4hvzRgFyv8Tpn7MPn5Tqs
6IG0UfMhJH/l1cZMiRiUuNC1rM3+q6aoqHUkIPz0O5YpdqekIsFWExOrqRjajO71aYQ+Ef7mR/ZJ
uuyFnsIKb+CvO3aM/P6Vty7KqCxFNrkpdkwpylHzRHk2YSoBtDxGAEF94B4AE8LwlaKJY2WZSJGY
VtZ+keqKjeOgGWAfDk/wBuk/n7zVhCu8cffAKOsYrWd6CUFPVhpGIvvrl2IFRX9IwF6LIXVXrkVZ
GjJcJk+w2SxetdaGYmVQlXLZp5kaxFrj/B/U/idnusvxMhec9gsAQ/s16/6/0gXldIOh727a/fQ1
pisuzC/7Ai6pILkTtGciJPn5kTJG1Sw8nephZj3z2G4U22gBf+xtakIi4ji2G/3GQXWwWUjlo99Y
TqNUKLo7BDwg2emZVZ9sHnb90rFu9gBtZluJQx7xumUBH9F9/ZDg6rKeZkArx+Urp08iSiEmE3Za
OB+v3EVTAcbjdbCm85goRCGG2f3r7jWuotJKqSnZR0iA21PDAHSqMzuJNECvsPcnw9fLca/c3nH0
Gp85ZGYDOBpFEIJ/kd61qtLUUTDbXf7b3blFqSBnt3j+H2k7wlr5GQFJ+aRRpN6pU6ef7Kh4hun2
gwO0I6hVyt1ktdcidDTNolEIDZgs7z7km8+gzxU4xUoVkuWdKlYDPnO1xbKG07t7OWsNM3Q+tLLW
Ri+ufNsfMccPzJIcH2jT9s9A/vLtZ1i5vcsRPJ58rgqYjX78QB6r2rxmgv0KWcSit8iPyVB/SAGe
5eukizIOh9c68wrZCpYuquL4EaC+Re2gj00BNrVjX4YajNchdSYUmaxD/QVLoofpJNe7LK9b8UHl
SyMOdO3HpO5m9zCpGg8/DBkaV4sCGgWcZlVgTeXaOWKT1UPhE1rPfJXyLc1dxF0iHagiDYt+clhp
fz+l5smt3eIuPLh58z+h3PuZrrQVtTT9wKysDLbv1ejPZuqvA+k2QfHzNTjYz4711GJh+VFsE1TL
bKYgZgJGYHoEoF8oPReoAPcKLhMWzrsxO4W/OjIMVglMvIC4ykMePOEoPQMhve/nbrlSjQxHOQqb
9NvmNKw7YmFtkoAsAuFeddS2FdxOYVXmeVsNjo9FWq71Za+OSjQIzXVf7yS3bMeeBwpYbsPqSFcr
szQeg3JtHsVbU7OKM3GqdgbzhnmoLb/QCOhNKG/ZnhckSQzf+oGZZ/Ia5ND8PKdI8yvqvhApLdWo
PoGAnW3SuCREwSmKh8ttntrpc+nnbgI0CVz0gQfIAdGrXmB4XQ9WIL/4TeK+XIWoJ1rqPzslFK0u
j1UA2UkQpr/YLtWzbfpkowOuQxgjqKXHMEKbbperH5OpypTtu0NhUqUfAwV0cvEGy2Ac5Nhu9ABb
0d9hR9q3GZ79CxehZgJt+z2r/GEO/dE16DmUxN8lDEwl/99jNhF0HA2EVYogrl+Xnkk4Ofjg+kLD
E3TC0q/joVu881sBr5KoVaRHL56PNFXrPaCrquQhvNLHzXLc1AUposEi9BaWCrDBlfcX8tNP+Xp6
DLP9paKrZu2oi/fiP1yrnAFfGCrFB+Uu5N261yhiBcECFjXHPGUHPYO5yObJ3vPizuxb1ExTCKP+
hXb7tVPUFce8htNtQT5kpaw1sFzkGzyA5B5f3HeYv9Zc7ewyNkRiPNh+u9GQvFxbsJD9/MhrG+dL
7g7JQrRV/FM6A9Wsy5R7r1xpUCfq+clpoeiHzcKWsk3r/u6NHvsbfY7Ozy39+m0q1tlyYWzPEQbj
aDzSTOn4nNYVrcFnCkuhJ9Nr/NHnRP3R3S+u00QTzwfGty8OJawjFrqi2v3w0+Xx3nQYO8it8IaC
SD6SfB+AIifCZ/aV0TJwqgzsyiSB0FDoX45y70+1GpCS6lMrS/ehCLNhbRc0yRG9Cwy23fXB8XR3
gAz5wraHcTE9qKrkU8yUf8N4DC+PA6/nRY5/Mo68ef8C8ccicm3O+kB6bzc6UUWKKkGKMY5hNhwY
7DY1BzwcFH0P7KaYfClB12jymZKc3YWvwWIcwEEhMV3u/dKxH9mBPbicaZlrjejBBNcHsyWGRJXL
rBUR96fg6eAfdYK8xEo4p+btbDFm72Rywd57RZmI5EKEmojAwIDnqPnyfJGCOcg2tUHX0zGql8Rw
PxLP8YI6+UkEbs+7apQyMgVtEDMW+0t0Ib2eWc9nIXn+gAzrrx0YoMhn3RbkJsgOlBb7pxkRsdww
/rRfw1I46XZlfMDuqudGka+NCNIzD6E8hUW0xm/Z4pdBgwljas2FTVKGOe74DH/yBJTQBE+HNUON
JKiqnU0d+81FhtKoKIZxGK4V+vb75gt//YilIHNgt1nNxadviq+5++Q6QZaeCiEnAKwRtfbu17QK
7ZasOjLne5iDYkcfKuAdAWCOCTAIiDE3cnfnJhlDz/+ElFK7nemTdSKC40tXl/Tz70U6J7CGa2YV
bQTb1vD7ZtQU3wNB0LP7XBe13FdU29EGvfQYSkcRp1OcTB5F0erZu/MhE4n90JWqjOffIvL6rEKN
kIQq1RB7o42gxFbAWCXuckbd8FkryAHkofwfJbcPxbe2rJp75Pm815+sBE9OluRA9kFW0TqtjTJ7
74CRcGEugvg1VPnbmtnYdVm1Ta5f8r/RvYW4ESI9NoLn5ZOgA9Ah54Ez+g8mls+B8SBJajntRuzv
n4b1Vft2EJy2EQSRUi6u+8weGJW31Dlw1v5oKmxWx8UJ16hgdvkI1MUyZY6+tV72CkzXwaFl3vlO
BXgTAp+CDGLkby7elAV+ePv/i0TbMx7u6L/oWwdJH/Wt/4iWUew/f7HOsz4dY43/f4kzsSD+8GLk
0IzWE6dMb9vE4E9zCyYVyZDtLJgUSAVNExsYc9jZpkckQp4cWY/+3niQn+9Bkhn7/fC9u0/IW4aG
r/LA02B1XYrOXEljg8feQ9YjsAxzaSvMxtSCJbd4pnPiLY7OCVWzfUvjEY0ZYv6vpKCFQbzdhZIP
XQXe/dhz291dzxL67eRwkXkUIi1NKgLu9LGJLUels3VN0RhNE3/h/UzDWjs2KXNzGP4hk3ivkLtX
UGBSMSpBbTUpom+7/4DFfqfw/iVZvpPQTryVIQ5KMNzSHZ11WfmCRzN4J9Ap4yfoJI9oGm63vj6t
h0YMsK7bBnxMKglOci2mv7NHMAhnfY+S2UT9zJ+ICOXU7/0fi3+XJYdwd75kjR8wfjjqHgPSSYhO
AGWLU2Fs21IHvPUeWaaFa58iHU0GFNoQnIBQIq7p+iKUAcDS6jNNFYZIHvjpWe36Y+hs0ARJ+Otq
SyYenlWXUgtKXWBEPmKUGl7pM+myGy8A07N+bfRTLUGyNqHn+tr7hVkUy3mRzncUgsZYwrk6etIJ
RyLZG6Vu1rNxKZuePzGn2dXqB6HqLVVfsQ4tngZbgzaa5Gf/1BWsORrLyu8WUD58ftUHjlwj6Kbm
VBiCV4IrDokz+5q7Dk/ZOMzY0oH1Ig5TBwcaNzreMW9gIi6fRCHecbZoq7x+xebYKluRvJf61s3K
3MPvMjh7//msrfqibsLtNijBNUUvcL4UGtsZLHK+1bd4ica023OZj4dHCn6nDiV0R9eiKYGOE+JD
EM4hU0Oin2jFHsN2abd/9wwci2lwZWqeJwvWVZumd+sWFFa4kddJPp8FfcvbjkNhEABGAQ8sfx2h
spQS041VbiqBUHixJhjB/uuIXFFYbepUz2PUO4/mt8HsirXCxW1IRc7HR+qq8rPAd0vvP8II3sX2
Ibgz6wKIOC/RN/415MN24pssEFFJ9Tz6fdN6CpY7sHOE4ZwLbzIpTiKYEukOPadVrylcGishl9Fe
s1bvpxOyPx+I/rSvE+UHI+/51Aju1lGMc7dmUC76wS1r9Qy5PgDhK5MnH2/3jVj09aua42wb3Tws
/NHcVAkGNfaphRsnRl2UgO6HBcZNBBkfaKMx4SNGpISKdhROq3w1KPSsQ4gcbSNF7iZ2suDjyDtF
/Q1YR5oQlXPvQaFmyAhIINslBzcx1AmZnBwqOzZxoA4UCslk8hWyvK54wlReCLB9L1oftEtw8I6P
uE0VwsN3wYiU4BSbh0i6/Xl9BAvlBScuHG3SdM/19xdp4fnN01KzWD2/zsLnGoXtHcgFTfOXPaUo
sKH6kMTGJLbcGyDsDns3D88JTdbXvc2erYNmokn2XgLAjavuNQXxjpt52kybh9t2yIyVMjLst5wr
Le2maUo2wbmqN6Xh3ILmbFH5j0rJUixvejM6TwtJI922p2IsSpCkNupyMDZMKoZSUA/rBWwqPs6o
3ABdf1ely6Q10hBvUcNhtOxxK6exnS6DeK0cm5yzm6rOQ+nZDTH6oBeWQYnODcHvPQCmJEAkjSry
SBoIYb6SOigfTpgAKBHrj4SyPxRD6IGE06+70GG2uUlhCHLJU/ZzKagxmxFFM1kMtFRRQkBVaXU5
szKZ85521R6LHnGZl92zQmM0yZdNhBOiJKqHnAtPUE3NwGLigUmfaahjvsnSTDFdoNhTF8N5Ub86
7JOAqez9NrbX5Z6LDZCfQ/ZYR8wjztqhiyr7kYHKxN/YraPkm6rgVLAifJVo9rFCtIxTNgMBPKGH
dCOWHw7BeUZ7HqgsCxt+6AdRomKgjvSN3Y0WY8pPcfJZt1H0c7N8rLRjnRjfX6EgtgutmBPlQi09
5S9vkJhUcDMlwK2FkqDXqXe2FbDX6MK+aBs0R23zMBfzjzZByh5IIlllwNJBcOMSIuYkDyZR9SF5
T2M/hMVSQZK+mVSiEYqOIcQJFeEA4I8UwlZnqqtvypuavHzcFbjkuIiLMAlIzky9rsBHKgCIR+iF
BB1uM0xlJHNyBLmRAPcEGjBUR9ClAnYhgJ+WFdnqu9VndPxUCZzR677gdhaQUOG8aBa4wktiz/Tn
jsv0kSgeOoSymiwCvWUw5UVglsObuqywec/TmiKZSjx2Vu+dxgHPaWg0xuflPAap1982Ef1O+R7G
EhsihNzfgpv7RqLgR0AxfnOtKVNBL2rCzaeyJTHLxy5TVxSrZwAptGQmUWTdciDI677ERP6s+E8A
GpIUsCB+QA4s3qKtObQz+SwDo4FYj3ZRE0BsKwIKd7SE/fkFPwkEeXlxIsgVDwxwtlGWxpbFrUvh
jbs0onFRJAYKZibR5FQtUO2Fvo/bPIgl/GOWaU8UnSE8v6bRMlPD8AAM/EwqgJuRGCLrCukX3miY
zS8oM16xZqXCW561xG4feCnwrCy8yNkau+bLajEOb8q5r3PNYVvo5QbOWunxHe4CzI1hWIFvPvIM
93GLDTdCeS8A0UK7PhPQu75IM/DJU0s4wQECcccsem2mdL3yI3IJlWY0I6m5RU8pvDIpHkDsj4ZC
LEabu8NAsHgzL/6qz+tIE+/f5CYZ6VcZU8fltz277y7vNvL0U6KQXRUlotkosZ64tWNKZNpEyJw2
fg+3afjD8rCZWIqlM7X5Dr17+m62a8m5fECE8DnOCLQCXsCd5kr7AYRaHoAFZoBnyMeEnx5ckRS/
W5m4h6h+28BIbXprGqgo17UrShLwEGBS6mcMju4AAx7TrokWaA1DJ8GSXIWTIZPudSJYVoyVx2pR
NjqI3YPRLvyumdq2GGhXFSnH42M7Vbr2fUsS0TTYvB42DeoCEWG60D7d7ihv5GRkXJRrIPaUhuby
wUQ1qFQnQ7XlZA0LHJB2Mi4cz6BEp19UYOc5TYzrSaHu3gwWDFlFahfXZrUah0CS6HCo1ZkVhQjx
KQ4TOKznG/W6mq5YyIWmlak6sdvY/u7PAGpBNhyvN9PfOubtRBbHHFXrRBiNsBPCMchxsf8im2lb
wKp+FevA1TCC/lNL4FAgHdbccAn+5S4/RtfKJoFQdGX1yetnlqBPmPAvmgoRFu8Q36OzR5S1elMb
L15bX3/O3GLA05Lx37A92VMssBf8XOvsdvKAbVp+YaUIli8LZGE5HqA+MPDE1mHtY5JhlVBDoTzC
ZENN7qcTIiGiP/PrHXLFaHYLCXM8ii/0MKOxw2kdwTTxNYt/lCnipXYz0wGftM6KkLMya6GxBkSc
ElNe5XPjItXcGObI5tHfcpryQcs6EBjG1IN72AcpJbRgMLy/nMP+1EvJ+egVi0EjUrZHy233fcG9
bVUSygpha/NzWSLVBYZg1EAG60AK59LY4to75orT/uu4DEe77O0Qm98fdBboWcOA0kiTs254hGW/
N2XoT7u0jJ9JzzvYl46njhePAZBZa4ldsEvJtltbiB6maw+8BvSgq4OqnS682Y47Oj0/m6y/PM1R
2f6uUTdCEOXHE9U6t+FTGPGbOYJqXUsFAaU+sH3ab38LtbnmIY7XFUKzIBFBPlkJTd1YnaSPy0bL
KDuSuqNhxyRcDQGaj0gK/lPGJ7jt/CvIqhxkaA9myGrZiLiRgkezaU/3U1u7aOX2WFP/o9znF2qQ
52enzmNtYjdiCdaBgeVymQmVhF3ndZzeSfY6w+Ifxt5B3CXN3KfeZCYleg6HGBKVVgVBCAX3O2By
36A3IrXJyHGtlMNj73L8hKVrq7rt7+L1Y9qOgt8NlO2V4yJD3YHr7lZtwfnNHMTLjHpDB6xtEGB9
A96BMivARF3uATMGfXe/ihLcJbOGn1FFnHvWXouAxFdYDEN/3DDF1Ht2eOgFOPOzWhV5rPe6IRrO
qJ1TwJOCueV5D+GnsZqkAetJO9MGJf1JAuJMQz/59Kvej8w70TiC8ph88BDjdZk6K6J5YBz/qmls
+NbLgXQPAbmMC/G4lZIaLB9ieQ8unDc14pLhscknRh7d/rJQ7Mr50k31diN7zGeAuaLVy+lUkQS0
VamLUU3qHwM5d+W2vMAESkrX+Iqg9/sHy+7YVOtJnCBe+NqkC5lgSJHuOHzLCDkveLVjBihuP4aN
AOWAfxa9HmWIC5UFkbpPZj0EJYOnMTFtvW8riGj92QTjtM+UqEZuPzKU0D8fqYUSU1uH9o2dQ1UO
uOP9w8a/9KibqoMmD3nTo+lNmen6TAyTirsEXy1eBcp/yjMg37ajMCP4hYS2Q7/9uBCEBPw9HGeM
lkvOeYcamqujDMsQk7u0jWF5kXlyiTDYHOvnxJQjWutqNFWhf16PngwBcxPirq2lg+HqlEz5ZxJ0
ihk1yONSWeVMSOtuLy+pqcBfsQO0XsOMtSFJq7Wiv9JA/Wz0V7A6zd08VE56yDbzklrKc7leKafC
rnfxLYmBWipY9ho25B1qHSlulBSS7XBPAUEzxRbPkJIhkoXsBZWRd9ZPXnKR3y+huJBzn59duFd1
IdveNWr9S4aLCIe/qvIC0JIT3e2wgH3/gajHAvb3kQQKbDH8GXCg6EB1sExBMEm1U3K8Gksiee7a
620jyxMm3CcI6yly1ssLvD9JzOvEcEDVBP82DhJR4aprsCp6K2n0IVafOhZCEEPV7RYnDnkd/SIR
vLcjZ3v1ndYToEffJNJeDrwRO9XPsV8/NeLQCkGrbf0nTt4bZh2IseKzi3w3IFb9X31dM4o5g2cx
MunbftjAsg4i6Ey7lvS2tDz5X8/rplx1ExH5m9Er2jgWQe0beb5t42vCZ3hd2kIswLNOgjnKa6Lo
TqsEBKqDCrQLl9SLvwaN/YBkwWSV5IMIixnN6CaESawPLBEkakoZxLczOpG/V/Q8cbVLaWLgcLFE
bjZuy5sXyifPSgSISKCPnzjSUs1u1Epa7Qgxo2xQU5tIkdpI3sacpsR6vh7JXmNXUwLX7NsZCabk
OnowUl6Z3c/3FqkfFIEmfekuKOLK/Jti1vFre60fXmn6V8pHJlJrUKmpDyQw5DcuqytUN6nNMB2u
zcVXylOFdPHzpD/oaDtcx4Jm+T203rXWMJ6xBaaXZwbz0CToLT9EXQTaK6fOrhHPvFyA97cCNBg+
xXCdtZlD0M1G6nMq7aoPDk5IN2Xxh8nLGSKVrvQARnK0n/+kL2F2vkbUZjgLs7EUlNoz/OaWYq6y
dl7CD02ZMVQ7Omj+qxHAUZ149ZEBGVasQJ6IorHJMBHNf7Le10b+liuRPkzF0P1CsEgHYEeehj5m
L+jypJXCasqtp++QmSE2XKASMHDCXPSEZj+M+9Zb1uAQT+HcCK88Ak/VZi3YpT6YDBmBq12vIAUA
G3ldDWTb/iLeEZts9t7f3BgEMk0oIst+hWm4ZSgcYi49pfi5AuUFzpuStY7iEGUlqrjMrSBDROI1
US4SwmV4SyYLvT0V09U7F/ebKIqWniAH0xBRtTr/PSgDIqVZmnX3RsQQS9AIzmd73pFc8WgZ1P16
E5o2/JK170ozd4egculsQnz/usbODK+0+zuADUy0uX8QH6B1IpR4r7PgymDDSlrAgPPqaUQlUY4a
rbLrgcfiZRCP5PtpFpabvFOuIB8bqFTt4jwcsbOBngVpnkt3jS9tgg44X77ZpleiJ2MvIWDfdHL3
aowYy58ZOvZ2o46hEBmzHCj0x6I+SexCSusjYEmTRpeVeYZuf61opez9PlNC3iQNbQsx2Ishzf82
ed+M4nWThuJ94Kou6MIKkXU+1kBGnxQgi4KbAVFYeCMVLaaWUjQ0GFCIt0PE3a0vc0WAL1JI02NR
P9vZHk8EeSqQnhqOUxTgYRvUI6Jq782I888VuMUZ7BAQ+NVvBDQ4jI+JvfEquNXAqir6JeXNdWGv
N3gzvuzMoKgU7STdjjhXHeMsrEcYIjeGFW8Ja4mZtFy4jtU+jM3KMMQH4Bdl7ge2sXM9oUGTsUsg
MJ6I9YLVjOazGUASbvjrXaHpctDtRnO2r683JZavZFtBHnh5Sb5E9Hf4QO68iTWMVTmRau7jw3J2
qjyDlef5DeQ0ATxyTy4qa2PLFTyMnSVgIsMpFYzkOF2t3tqtLpcS/ZNfkHPGW+Lc1Suwln56rOwx
SpuzIRCtTTR8ZPwT1v7+2+ft9MVfBkNeiM1ZFqTSbeHpnq4l2aSr+V4DMd6x7OaBeSKhkT0Aay8v
+Tn18n7FPhfgUyDmDD+Hg+9Tb0uykVhLSPGiwCP3XCe35Xr+sXQbt7Z9BiqtyRGEMLxn7TzWD0oO
DcSKskhMUV/a6W4bPvnbY4GMy6IXIaNVpFD0vElSB7zrTlq7OS6ZgM9Miiiieh7vMlzE4c8cX/wA
2b1wHD17n9mJIgjE+w+VkZqwrqm7yVjbHC+YNUDJ/FN75ZfQZkFX3k4U44zThe4PzqJDohLecgGI
T2risJqVD8uSd0XEGiv9saC0GzMAtHin29knOy8OcJn0O1hW1eCwxc/fIbNYVcpKqqhf8auXlMHu
MD0XHHa0eWVCWLf6vcwyxMjhGFbDGxCCQvVMuskazn7A4vyKAopYxCeJVANqxlebwPhRKVVsQjXr
8QfSXNJa0PaL3cRTAfDcKpaevyM/AhtjAvM6M1E4iQFyyRMtXiZseavoon5+iR4Ji74JyqJeJywx
U9Zsv2WOUBlQcJusUfepvkAEGbFwvtEyIj8y8COU5A0TCTGiizMHxtvaK6f3JMI/Bl2W0OHWKbQQ
H3S807LHepdsuWS4cjCpikU/f/oiYFW43g0agXn5qg/c7plqfjst72D2yNrM25qlj80zh9EDpYVF
wC28GVd+W61lUj0Zufjr/7xojAR51YS2d3K7t9OT9j2T+HNbe7yR5F5KqgQ09OS9sc7YpyZFse+g
a0zBFqcQxtq+iJIiMFXKaspzcN2x6Q6rrfKikCDJBlG0HGGoOKAlhXU8s3NN9y7jVx//QRYYfBhU
i57ZWkh7rGHi/jyeeIj/yCutU69w9/QAdd5abbpzKJ3Inr/oq3HazMPy6/I0TDeRbs4derJR5qAe
1jReB19hGvuUBT/CYtN7sTvnawAiLqnGxmi8hZFmjFz9bP1zbTMYSm+SyLBy5LzCoIF+lHBkw/Ap
LjMNabBYEBMhJwIz63KR34/ZZx6id66lQA0jkPIWCDwR/N58kGvIzBg4Wlm46fibCVziwAjEp4oC
LYE40XiKp/jwsgJB45+rGOQ76X4pWOKa3c2lI3B2zQF+J0eAJvcpqC66U9P1xbuWB/E7xK1zCvmU
Ne8Mo2TW0XFKrubU4UHnsWzn6+XaV89MWBVA/siypC1HLT8qXvZnWlWyXVtYTtrSaCE7foxqd3IK
Kc1nYIGUt7QpwQEeEDz/i3brCZuEXqTQnSfBKIvbnJD4vUiIYLhzBSDbn2TYG+rXIFOcOkmz0eph
fgbpjn/mXLo4XlL1aBAlRh9P9Fh+KI7b/EL602VDNRkJ0s0JC5qJYufm72ud+QE48gnuBjbRUDMI
eLtQQiNIIfn7wozOXEAUb7GliytvgKM4e/myw1qf6Z5dwXnjDq3D7eqa9xvY4TRKc5YwDrNNMd7e
EOx6MIl8tE4TAVLKALnbL9rMqJLIzroNt2hTykNONbTPwKCreQaVrG+0r97P0gDL7Gzdt8Eblqy/
g+1nYvWqV1GpzQB0od0XtlHUN4S2cTpUnUZUsfhHy8EloBiyHRGyxEhO5B2ZTFNoVU6PUPN8M4a1
sZoovwV1wMwzAImZftqsski7nCLmMzhauqrX7+zupS/DMWhJBULNYhUqrOFTG+/7X5TOYnqSLosc
lmh0ENPKxzQWCCEU88lKF5K4+s+9g/8AH8hyIajgJQVZI/69sihDldKNFS58z71/oXZogomjxyia
or+asdYYf3KT6/mPXUSB+lYUZtehwjT3/fwzKSEgcyE6CPRkh5kg4YCK7aFs6LAcVyWcGBguNPQC
6jzCqc3cPsDLf7KIkc0mmpasV4Tqbm3X+HHpvaHffmDJdlsRLv4WMMJSUq9yjqx4T56CtAS0qbWi
hY+auPXqYf7h4x6506BYqgKfsuoslvE+05NFJEUQ3om7oEjSnaUlxFwTovXtm7ngD9SllZERqZEa
kVHQTyGjQ2ctXl7HRn2VsIeloCA0U2QB2Mw0zxr0OkNE23HfD4joAB1IgfgIcPRqbEB6DgTtXwd1
y4gKCE3TFLXqkPsbma7xH2waeEnsruFsvuohF6wIp8sVqdIiP5dRnPvKXG0wogtsdcv0Qn9xn458
hMCnd4LEAp66PGieXKeCoiOEiC9L5wtPq9dfWz4jjI/eiCehVMbiIoqAloSbzhJ2SSItPsgpjEoe
Rt4dJFNTNQPJdcyqM85KW4xGT789FzbhQp42hegKZreSOJl7bWCXubeXZA98UroLr/SSfKfcF5Fk
UuB9dMwnxlPC0FCnr8qcBF1l7Mb53tZsz7pyfooZN+uT+byFr6hjpFp8E82zEzlUd6dA3lTPt393
4FGlyfhSNlTXRx0VHEEZ8rx7PcI+bsW1JGAP6pBmMryDh7FSEDDYyyXxtUEz0bZTccvZpqh7a+rr
lULSOtTPqJHE2e7/GTK1gGzduTJvzQmXQvd3DgKcIxz5U4WhH3r9Cd3AaifrvqcmgIdbmgonlLol
5QbSaVY0sNc0tlXD29HQJulTWWz26i6QVsYAtJNqG8A4aSmNlzeGbeA35IZJzzDVD8/4cEpmmAAd
co80f0TsUXDy6xim4ZHC8CnCtqaYZv/cRR0utgzP9BxMfKNq2obqfOLnW+ab2XLl+BfMSAFP+rAB
mKbEjftx/zV5usXhUCMPD9jmQxx37TOY2F253mV/mUbBZZ9INLF9qxSB4COessq+BUQeHA3gquOm
nQktIeRH3IlSfitrdnmRoy8EkF94Eoflxynx7znjR5NlVf2tqPieiVNxMSxlo/9T+36LTwCc6ssu
E2g8dQv6QDxbV2cUWxYbnfIxO5iU3b57A+jpx5RVF0uc89zzYJGOwVZ6MUWJKQQ+pBRaxohI14ZO
U1RLyyBQsmEJwcSmGI2UVGwARxuMD3UzGQ7vDVdsS6chPM2KyFwcdwCH2e/l6HXj7VCmZv/O5fHA
KpG8kmllvN/i/2D7o6us5TVUp1d5WAvPZ8SzWHLM2icEsH5nR3+eYd/+YKPXdzaW9ZMzxi0W8XT2
OXWRzg5mAZAx8OzLqGYnRTfxY4y0eKgNqDxABzJkiRwcVhDihfo0YqXGSjvhf3MYdTNfSguLTY+C
8ZfD+cAjGEoVzwwNen3oQM33xvRfPnt/rgdTgyWexh3aRgTaMvgx0oZ0+H2wuFTOy+66h3pVz78/
LM4KBG7K0ozSkq5EEtYZzLfjlWyCJQ8ajYYscTcYRmYWn1PqgJf0E+9PN+PF9yvd58mekBRpk5ud
NDbX4jbTKf5rpmpDHV+6FKhLrBxDLoZhlaq3gfqrdHUrkkPVHEsBx100TxdU1dTYmpyJKG/G3S4Z
9bkKBcbnf/OZEMCm3YS0IbuSaHDMGzFNYmm5pg/B6xzo/a/tQypFPwLYxq7qTtKSrb+Gb3TSv4o1
C67i9JT+hAVuVTCA6DD9XMKQTLYpkLkbdIKXCNchu0+Pq/RtIbd+OWqwe+s99XdMLVz/apsQX2bv
RfLRnRNP8GE3ErSxcdClXNmASuvFUQ/DDlugafeK5brijvPp1kNfFqvxyDQF1kU2vWRdtQIiApOy
I9mOD4h5vmf++VdH+2ZiwhITGIuXXBqGmkQc2JlNXJLaJi1cOu/Vv9CJfTLEurzlS3aUvpEIRAcx
QIR1AcZSnm+RzICQ2L+Zp6TO/SaBEYiML/j42QNHxApO6b1y22st7XJFF3HSt2LEe1RkL9KlwUUD
3uRlnDF4y1oyoP7mUpbKYUJy2mZ0K5/kDfxg4ymM+Hba+0+IltkjvrHfzVaUipdLgJeofeUwJ50W
3S9pBbkvCLlxbVhtbgpT0L6437bwPy64GbrV4UgN31MysoZcj2bfqSHdQFx33ayMdS79Qt+d8Vao
e/OP1aanX7dIzNhgZ19EkPDqrxUyQ0oinfF5HmAq3OUcXrw96Nmw31x6IXfn4b252sYQMjqq9cg5
d5OFpo0kecqM9O7MNsPP3cw2wt8E4KNjowHkDfuXGAT7Rd50GiwAMWqOI8dBFSOiqgPzIShh2oJl
v00FxosV+lZhG3x46nSRJ5oPsrIFj3cYCEe8tzmSqI5la2vY+UDZUmi6s9qD7FSCZ3Vu73L792kr
TkWOAHYmVgPjKwa3G6Z+CHtpVGJV5VkkBqduGk8YXn4ecHKytg4DBPXS1FsBeqcmGSWZ8di9MbJu
rmxD88yCK04fTgeZQh/ojj0tb5nrmvQL4i6EbaJUs8OLTDN4BzuyX3IhX3M816siO6hcAqjG3DbF
KVOSQQ6RsxJGKqogvhIfrJ9+R3/b8rqJfaqsxRsLKzc8tSPArju4xncEXIni7gj/D5Chg9kGZ22S
r/egTRpjB2ln5SkpojcY3JR8/QMcbuDuPdidYwJT8aUqzHPjaXIRhf7lfNDcBD03rfpuuhA6SVce
gZDnjlsSKh6E3CrKqb4tLojczkp6tqgzt7RSLFvNdfZBgFUM+Yu359MVKPc5ZQH/d5VnoQcvNqrq
lHr1lB4D9H/nD7mEjUmCqEAWR8T/FPiGKkn5gw1qKpfwzmyRkQzVXTW8QA53/e0QDSSb6JP1B1PU
DFLP8mL+cMT9yEeUqSXxUGncBwPim+tvYOXx7MVNfbUzro86ddNmg3IwSboi/11+HzrN+qKt1aZG
9iAVoRxEpqJc89PK2AmurbNFzAiw3EFRLVXPXsYomrb+pl4FDSSQwMBSLwtmOSkAPe+HU4bPO8Ct
dlvqG17TbPh93QIjSsDTwAahWSfKrnrp9GXVxgNRUOzVJBYa3l59FaPqmSplGN/88rvQKd8XtO82
ijdPg3iwYPhP36hheFL+zDmaSTgGBkU0dR/+xPEmMB905Rm2YqX2p7Q56NTasgjVd/6vB6rrf4EZ
GKmHVM3mCMjsrAAeZg6uOZUzxa0J+SaL4goeYavSYgmsTuG8MyBWYSHrLl6xpju+d/WDhy6vFGv1
swwh8ESLo0lsTcrMJAcLki+hKGE0DCb9MnF0rhNfv8KDOsRx23pzRVkwUal64qEsi0FCypu+5YcO
PZlYSMn1kl4quXmbgir3fE2E7tUqe84K1Cao1CGWH3Dr178BSzlBtTZsqsbLnKfwST6DyqlgRb6v
d07XO0tTXkbfmmreRARm5ij2JsTSw+8u+mdizsZFZBwfEZfelvUjeX2coz38CvTDVvZ81+ZLX3yN
7D1PiO2dLycO8EfdZmbY3Iu6YBPfqK44dt77Bz18oDvUlJkfZP05AilVgg2WjKnTJWf5RQVAzySZ
Gti88TPb/o1MOSuNxYZqz/1Y8jdCPzQFPNQ5pZbTTkgr/IZz8PNmFM4ZbATLMjTjk1EBTebew/eR
Pd1Jru+crmOh/+TGHxElhjOGLpP4vrlT94Yaahr3ao7Gp2uRAWQqrVH8oulDLotS9TQo1qJwBpVP
uaR/Wc0JF47H7UoXt7uhPBJgPadhgyEPXCtiDbBczYH05XN7yLQkcVqN+67FuZ+Q0orYcqSEPi/H
FE1E3h+m9efn1fyPj0Xl4u7ZJFAqKmuU2135Olv5EhoC0gC2u9NIFhyKmJ6uliGew8k0Jet3FsQv
NsyOM7bykJtMRt3391UBmangkKaT59Blp3Ix0AO3TwX8OrGdl6s992tMr8g6mxCwZfEmMeV6KKVM
YBGMYnNjl5Gwp0cxbCJO8uXcSzLV67gK09msJGBF4qRuAiwz5G0/jkcjBDjzqHgT67S5qJ3AZHNf
i5r3yNv4uaTeq7dR1b1WbuzWfMCW/wJHaWyDAmEheItFn0S27zWnnIRKhaDduADPh4WgINW+BJdh
Ig9rOi5ip8FqttibufhxMUKw2HxYw1Tt3hVh2iiYhEGTnPgFl4x1xryjVvh8J5Ozbx589H0prt7V
tzg6zKgcYLTPU0uE5UH5q1m4ycutxeGJ6URlI5hXWLrq5zbRWtZOlNOcApCLez+Z9j04cdHFV0T8
g9pfMHdWkUdiaD3Vv6FjCo9Dwo5/kXhyXAHJnYTk8JI/Dxn2QQjpXlV6Zid8MFZwdyyW6bc0oOOL
FzJ5l0gj7BK/49OLgDx8sCp3Iq+399wklIo3bdgM5cuJn9w/X3OlvAr5BuNOZJusCKdgiBb/N4ER
TmPXAGAC89cP8ckiq9uEoKiLyMxkh9F8ciEfxkrc5sjlpfOtREjYQkLTxFS3wbJqaueRmoadQkH4
68tcDWPBrTD1lJhLm3AU0Zlg2/5GRA3NaRWPekDfibbwXKTI11bFUX33FAIKNBLClftUuAv0/atY
OtitIlPZgwMFnyYj6LpG4jvr6lnC/5W3E5DoSryiD1vXM7QKrI2H9QnGg+3Y2tRAL2D7ZM8QfMUu
7+JLflVk3vmb+lxBH6VGdVorb5WroIpkgTCiZeEfz4XYPBng2ogR9ymjNQdaVBk8CxsWNSWnzN0O
7vob1XA9l3vXv1xCP2IS9hh+k1+KuJ996+eEhrMl23cfF+jey0flQ835K456tQnbn2LtUQtwIvmL
czP+mArTGTew1y1Oy5MPdLmFHbE0zKtcjSvF6mdmr802UoKlV6OEwdAJHYEuUskZOhMMGPwoMXTD
gBLkwKPSQJ3z9RtCTiSyW43WvMK+24GcV7ZiwapTrnUcDaXR7d0nVAiZBuVMALhy6kvU+Yf9uGx4
NrBCoczZmPmmRdXxBjR7sRtx683/RrjiZ5AMHqH8zOa8p5c5eRyYu/Raz4ePX7qt6tc4cUfTg+gC
QjDmnWkiYH3vytvfhmDamgAKTcueaZOqRW1K61xcilTz7oiaTm/vacJI9bWL33piAwdDo5FkOuha
TJfjNuA2FLstcZ1RytbzqtcMFOQJM1doraxBL6PFtsZ2Tru732NOha1UzljyhdvnmTkAUenjLcUb
TJEjxLpK/E083qA3yPBLZ1FoyuXlxk+7GCpLtGh7r09/Xnv9ls/jj4q4475+cQCRJxxf9UNUZoV4
4psgk5G9ahOYtI4/iZE1A5HeV1iPF+YvzG4znut+lhBKxedoqoj6EiDDBidREt/hs8X/LIUDgO1J
Gx7Dv8DfYCb5wOzUAafxxtm6HqoZN7NBib3zxwcPxJK8SDVsyfHJbcoxcj5qZ83eNMZEPWv0UM7n
y8SmUMO7UGSA6AUjkvcEhwsHLP3bcd+bJWChMlut7/2MqrasVS+kgjuC5zozzizQF93loFBg6Zq8
HYxCB11AJHjgHtfoxnDtDEmPEFIntNztuMeu/KuMUGz+mWD0jFHsSKespjuC3zL5y5U/GKxxqunj
qL8iIkRlmu0hqJL1H5jx0PxOcgJq2IWajMuZeHMsYBZEYRcMQlpn6AEmJFFAcZcdIju155i1RLxm
5X6pjNkt+PjOVjFxA4BxoY2xFbYnDo6vmI45q7J9+XHr0d9pa8XWPhCpF9uBqk99hfjsprOUh2L8
k06Fs2EAXgHTsC4w57GxWJPaLwc07Fb6O1P54JBCjGwrLW1I7QC3H9a1fnfb7WgCTpT1fR3E0lgF
a8K7GQGsJeHnfq9wrwn0SgezSCvzGliWL/uvDqVfqZfMDww87+L602duZhOuwEcO8ZHRPILBV8N2
N8ERLoB9HsAISbYnGUil3cJVBxVKoCUFR7l+J+mZlBwUWCKstYuWzMO3nRwhSv/3THpk5si1S9YO
x86SGNC12mpT1BdLd8r2ZWrPN2NM9vfxjYwyXepTx1ApKvCsxdp9ss+54mywPl8d8ZfrDS6tLkj7
3hm5NO5FZ2PjKjSuSGx+RRE3Spm+GfDk3btqC06O6MbBkKXzMRjpuOW+b5jMsKJRpkk78iMsXbNt
nS8uHl4g+ajAtZrIOCFiaV5p8GjpRU7qu88L6AMTvlwncHUCSR9ZWuoQN6cEkCfTJZUZqAG3fmGM
Tq//oeJmu1kM0yopUmeRqeExPi7omF6GAIjXVNY5R6OuIcJSheSVOfeVAX90HqzHrEwIUCVB10ig
jk9IAPRiapIH1QajJoVGetGaqIEUn+YmGW/dXnLl4q/PM0dh0ryR2t2EVExRNX5CC9Ii1eGSTxwj
4m30HBJb5WiWImLfagpc/yzn3GsOPk02atqikqfCpjSUDg/JObFkR2t5D23Gj/wLMPxdqsYSW3Nk
9G6DzMJBbukfIOfbBlK7bQWveh7yGjnbgH4sWfRko8Wm2qyb6xjX0dgwUxRkz8vcmu41xk6+1tTo
uHn7Jes70i/Dt0f9xR6HoY2X+Zzxm0lRC73I8YZblBccRKYY0b3VTTFdEWW7XIhSrDNj9G6Y5D0y
Ivn326B2UEF5AyVH7/Tse597RfrHZ/Mif9QWrURnuVx4SJXy2z/kyEDnnzq2ARuEH8dM0x1SYKI5
Y5sx4MvHFuDwSBPOcd228wqOj3I+eKrCcvn+u3KuYJYhiI2PgannKOnxoJg/LlmxxjCrfSpYZiHC
l1M99f58cEbmxiqT76uqYCnTfHzokJDqGFI3o6xeqVTjmNx1DvewHWg8T4nhEJTy54KjexYERdho
Vr3MFPG+PO0/IBuuH5uh4T1S5f/626bL1SCVZG+7ZglFnsXR48PkyjoD7ZkuHIEEQ1RNVxt73gW4
N/+vjwZq0Xd5U8F96BNYh+GdQ1aniyloLsBMgMA6zcZ0qjD2uyEu8yBBlquGVBWf4usojfiPUq3U
sVLl/2Yqfydx4as6HMmy5UQ7OxznG/KPqd8hZq52WDZ+C8iBFZx8qt/xLsvSd0zFFZhk4NfGZaUa
NhK9nN2rLFLFpTJ34VgK4C6+UvrDY5bVzu/+PiL/sTYVHZfQxyQTELep8mmDkSqJ4KuSReFgLaXh
NV7f1U2Ll50pvGCSWsOGlUabJzUgbtpuRLmpI4YmaCf7I75Nbph3fl2AmMJU8UpPoD6ThuYzEDz6
qcF8up/LpbESVI6Y5sdm6B4ctqSbgocHyHP28OaVYvYk17xAnJR7JggBpr0VgmRkKgeN8cJg9WxW
w3jX1FL8f/9XimFoes3fIDN4Vu9S4OBEBO4LBVmYqt53cGAeIOupKRjzVOkmR40OX6Xj+07ZaP5r
BwhVP0ZvWLwZhBxIlDx1g8Q7iHqqBA++Vku39j1xDMqvb/yva5MLXDs0luyWFjVzVHvxjXwr/TWT
v2nqrBrI7uvTDIgTE3/KLcFfd+O4XfLjgBUVtPr3h9+QKUBnhygVD16ypDpaW6rVgy+wHfF3Xyst
GngNVN19Bg6Z8k/WS2njnLDRjw0fawZwnz/MBipJF/Gm6vL6xOxWQnfMzMvpF7GoOuehTURBISDV
OKZyS/b/Cs3FeAzf8IH1ZIIBPk8jQro6wrULf6I8NVXk21WOqlbhykiaf0Fionf9WV4vPedfn3fv
qrNjBfVdnnzBAoSwgLWDkwX6meBMFX3ThFlaC65sHdfw6F45T9MXg9sXi1uBYuZfWIT40E+M4Rpt
rwS+SjUaBeqySoH4d2qikgJagA4p84+xRVmGVTW+a/2DEHBGYnhY4FgArNJliX3EA6PD32IzBCwF
g7wN7qozSCw1YKROvh5x1Kg5xsEVBoDJmKuQfgufGTuaxEHemY4y4U2D9+5paKCUBVuf/BvcIg5K
anIzhFnxbQfz3JndJBqMcDpBfaIjLT6sBpWtMJoun8dtYWkNq46bILGZn+eeWd5wnZ1sBZc94spb
DD0Lc8m7Km9mmhaCP9C3LC3sHVU5Vb09FrlbHwFQXb0Ix1NatFMHUCM3Xsy3zJwzCSO71lZIF8SN
m83pBmtNnvO0LJy0NvBwdfSdK8yQBdboRbDuaQeqJxXHr7N0IPGrZD4IVKwdMVpOdy2qr4ahOMDs
LvSTKINnRcVU2lcisA6qolbaI/dcRtNn94HkVcixyjevYyHUjMcciaQGiAewtcgzqcZogw2D9Lbg
KDaQPyYclFl34alaDN7p35EnQrBLdZHRVkYYtAIDDH/SZKkSSdI+e05qSFV2N07PnbX2Iz1q4TM3
zXyXBFTuEYI0YfxqYRk927JonFEnfUdHyW/K9nDR45ixeDdfoJ7X9rslohsBvugPqip8TEhuBov4
XEZC9vQcC5EkNsfg5C9z/VcpFvgtle3eSlm9QkG9B5IW9Mcp/NHC/GoiidaUffahbTBbvLKX81qW
50uJYDXALJGyxpmSR0XMJxMKQMk6ru2N1cti1ID94aWt1xNrZdF9QPkyEmaXNw7MxXHcbx0XWUHp
1kPuoFYWTeFmda3QnMLhmNz2RFfVd+a147U64vP5Fdcp9SbbKtQe27YzbvCTRvE3dpA4/D/hnMyB
E1HwvGOlalAP/RRTFnOa/ZwkhDYhnG/pWXmjdsTcydDs49nqxj0VfObIq+i4kXzW7dnPTMTIiNVB
ftx8U7Kfqw8f8tSpQI6xiX8htQbMcsGnNEqIhSfFHYTWvdjmWOibswnMYSlvdpIrPjWcoRFMcAQL
VbGuneQijhtZw2vMhCb6BP8JjEn2g2nUG9OrER1IzCMTiHGbzT3LSaImrkW02zKfk/IqlQADbYc4
QTb2flWqBZU0s6MZKJirCbbeZhVhc0DDXtd8fnVaoL9jt8qAVx4ipz0Qw/iG1CDJPkwMEjo8MsRC
NiDGqTLiZIBz3/qRewkbI4u2AFOc+gDbpZjz66343QI6FQlEa+fc4FoqYDAyEF73GJaiQR78mMwO
jYaTM9TJbTEYVJxZVykTXaOY9EbUZykvTpYNBqWYdrFMNeujtxj7VBbJ/zGU/zafCgR4wNC7bXdK
kK7XDolXmMY9fKAzKOtcDGtoYb2lxvbKMOQXJ0Et6+zAzyFSfECoPobKEgPCQYKW+C2M1iuRpNX0
VCf3O9e34y/intpXD3Z5Zwon4HEfIJVEN+3ehDxXUUfUISNCKFIfUUsa//e8FVZ3lv4DpZQNtx7V
vMAHF0DHIYvswDtGylWGbeB77Lm7yrloyTkJIy9ZSUlVgWiSZHTHdKGceRz77apTCEdg6O+KvCVp
FSzzICj21k6I2h+3MgxRfgbz8689opWifgnnAr1rerl12Vn4DnCSrqNrqJZ5QmxY/Roxg5ciPzVa
je6RYUgTd1nXtnSPcSdUIgTxDlaPJ8Ist0oi2k1NqpX3zynzOzFbb2tV7JAxQC3pM/TbTb+6YXCT
CIafMQQ4GmVDzzZeiWUDqJvKm7Hl0zZR8Ua9MArxLwaBw0BVLCe3hm6lVF+aVXR7irKvStTwgSpe
BvwsE7h/v62RHd/Q0CCLb65hrcYCXmRWc/U8l8mtRs3Elz/3p/aVTxmQURQFJf98B8gGilrqRqRP
fxKjJ/2uqkQhA9pM5RuXm7h4vR0EDbWY5jpeAjW8Q4NAQhJJLNTv6r2+FJUcdEjCgLeOujLX0N+K
0GUWRjTmU+oCuNbmVMalcrvdbTFOk6zPioQUrMO0XDYwL46+VWsIyoD0lH+NbX+IMYadZQgchvjy
frmeEflS+11X+xNhbqHrV7WDdxomGg+gLLuvuZodK5ebNR2QnMY7PdggzmKiQZOmg4NG4M1J2EDb
oMmSBtbJ5uvedainrAB9KTVr4iEHwl8exAzu9rorVAEEBE7BVfAMDJ78gLQRXWfsB61IxQBxdkQp
1qtT8bJ21iAN8wOoLqS5LC885Eq49CY1a7Vih5kQcfdWGbFfrIv4nAEDF37uon6IlSM8laGuyXko
LUNtBXdHXyh4aRlE/iOBCvdsvHDHqE5y+MD5942ut61cJ+AeckNvX4UixgJmpOmQma5ZaVgZGC9T
21UHsu1YSXx8D/k39miy6qNdPpJlKLBhskbs62gBiYrgW4PhvKEqAW6O0idH35A0VXcp7UFIHSwJ
V8HNazuRS8Zjo3/I7iaTSFg1N9K+4UkFCJQWpVAWQu3o7g9S6zidi4Oq2jLonz3RElHNBRVUZgD4
KUsb9KaI62/LKMm8q5LDoCds/YfC7ZRCLMqhGd0DvgW04Uof50uDy8q7qDsCzyMmDKgmjFxxERQ4
FJDq3zq27K89kX+yUbFYyjeRKDXQ1o8TtUx51KMEo4JOc9jl58ERszexZvl4rjaU8QP2vk2GMG2o
vFfFqPLMTIjkSxaN3KuhhTNU1G+Tn3jEyTSidZiC+ChMU/yRQT0WO7XDHb1e/2zo8MIeGQt0DQfM
w826U96AyFth2TAKW2aWWsZ976I3AKskU0FTAI5XbExA9RJzQ4By2DsxTlfwrMH89jbysSNLb5bA
MQRusS7DB1jnIeGg2KvZfTMETkwKt24Z5E/qrCayngUXzTu3RacgtugYXBvLOLC33XOBc9ps+Cm/
DLocNPWLqS8BNZJdsKcVyLlxcmLBbHhl8XBwbzPNkEh9z8Ihqqe1KUhcscJQPG5q9SKwGwLphCty
uZKDRjS1euvC4e2L02v9vosoMGo3LzB2l7tJiV8aLT5eFepHisjbtJI2XyhD42D9ARt23+DS5tyo
oEU5idhrPKW5GAvLMcKVzfyy7oUzhiux6ZBwyn08xfSrxZj4RS7mxyjplesGAXCdRAYfm3hWS9R5
825MiVlzmV8Qy5R2hqg9HF4U2+Ii940qZV6QLvjHcxhtsHKp6Sx87Jom032tgfal213JumcVq/XC
Bx+Aqnb2onL/r3YMXKnNxdq9obqmWSYs25uNshzjH1GbHA0D5ohEWkYvWitesT9UwlidGQn9aPQa
pupfVf4Z3cvWj4HH9hBXJHAZnMLjVjV73wK6avhUyzHXN1S0k2dnv7wJ++eL8RnJo3cmRHvut/+U
sbzt9OuJV3hzjrG4cuV5oiFiXf23PQvpdtsqLwSDzT8KTyOdyA2oii7O2yMTDYeGGVpehb96PibR
RsSITgwGby6vMv4TYSGaa+ANki7mx3g8Q1/oyAnG3c26QTn5BXf174CYLsRRh/heyJyoW6pxDdNX
zW/kZcFMlWFDcVq3w00PjptWsThnHHC8INLzI0TzYy1jU3mF+Pus/+pKOO9cCDtXKe4Txg3haiMq
74AL6j7krVKMtcaT/hnd+3+86LIuHIdgmK6x/8blYMJqCoPurra7rfNwEPH7ghnYJAMPhXO7uZN6
XWWoomYxnQwGCYHjhboPp9sE3khOk7gPlKPricWsXZztVUdACRUhOzoVVcrEwGvM69OWBrDeBEnG
4BVDjt/m1Qqb0vYMRn6ng3SaTBl0RPW5l8LZBVlDIcSxW4+NLvbj92V52l0kj1Fwj7MxVqwhj9Kj
OK0pPwS0Yuve4tc6o4NeB2nPNHCBn+telz8jWYuvVRCkytaGbM0tdNOuEyxs111JLbpOMWnMj+qg
I3DZmnP0ScyANZMqLgU7Tcmk6sdDqSFqF+Blud6R5JYMkyTb8Nw6D1C8HE+WKUPkpGiS4idnH2zU
vAf4GDnpCGcePepMOCpHvlBSE8AKZ08hzxZ+ZMNHjoj77j7GEHB784UHpbbH4jzvIiQmFI37NKWK
2JbllGN4aE+fKVMkGQOz1jAtZ/Y9TRzAS6SP3wobJgVgVUTSS/2G51VO0fOgNpr31XheDRqUBgOd
ozGg1lEUArI7xjZpBURNNwN8pZ4sTg/NfTqACndkCC65xrMJfMUwMHDiG6Ka4DHyZ4d2U6A1mFVa
lhBNcW7OdRNUwpg2AlTbJIIt0XWySKWIFFEKqwX2C4fx1+OpshAfZwRLqPwS6Dexiyj7bQyO/907
lB0wFPZnIZvj+RRWnXFhzBxDt69F2qUZN1pNvmgjk41aEkK62k15ptUlX+wIx01KYQvsUZFW8U69
BXu8KHwSYF4NmpIh14ff+i0/0fkQYkNFvPP9nNLkY1c/2XgLBTSEWIOTob63XKo8hCC9/4yr5LP1
1sA5VSxMXqyF9TS7zaZEpz3CzBmwJkZTCwR2vbyINkS2vTvgAupoDMb1yBVnt5SQttmel71BEvYI
WWkwQqxaSaKbMvOzZcRItObylmEQu1EbEqeldI7vCaPSZ1X87qywbM5NvD/EzRWimy2aPJuP5p/A
hQdnYkqusnqmV3slTMr+rgJY/wkjuAqJ2UdzRwYMaw1yrx5VwvhYJpUaNo3lw6aKQ9W4CFqVwhs6
TdoQ5R1SkmY7jBTqPEKU0/Sjp59futI0P7LFKGwbLOQNH+cWh3smyP4nO1NchL889pLFnc+usE7P
m9rKB4e+4L/CseBKf4WjwV/JMHpJORY41QcZot8TBGv9BmUP2jorGbPsKR9+sd4p9m+wzUocaLf4
3JH0FTiKfb/zwDi9Q2e+mWKMGKIqO2s+PSZNrnwSKy6dFlCtIofbUSLmEFp+YWZH76lsUlicmzRj
B9nBlCo9bdmkFVXIEsljAB9vigrjKE4ZfI+cFS3i4bklMjc8v0QsavYS/Uziw/COQwMcwg36kPiZ
EAVbDdsqIO0IzrrkDht6zM+BQcmBSAAk6yQWSm05B4TaWXiJB87WHC72fDx47tPwp5dd7Eo7Tsrs
ewHV6coTCVmQNqSdKkGK4HEDV6Vh6rc8IdEV/F3zsoqnNaQAo6dvrWSIgZb5xuZ8ylV0hBPRzemz
KK2f/CfkQQ74hdP8QBOAsmobllcewv8D+loZCVIvIv4MclBFlzr7nFLXNrkDrxQxrBsSORuThcHA
mUL3lCvXoP3nSby+VVmsPq1P6e9ZD3U+ObGIrig92CFEWoPARatlbVzk630aAzjS0in0k5KOOKLV
GLI1YMpjilAf8XnyIZ3GdErqGtgjYkxUgQxbVVl5DYSj1l0puiUskeLhhDtVGDT2Xr0HWe7HVEaB
Dtmdtu00OvOkryi0QF0iZBzb3a74/+NQM4KFY5mSlaKTeo7eACc2mlAda/dLnbRQ4oEZ11JntZ7l
oCRoW2GVzP3hp6s78eosHztuZYLQsyUg7dNactuzOzcQrEgos3SwgHPzz7U+yvR8D0nHtQZJK3FW
WeU4ZNxw8PU32uMc40LYotxufizLl1AwaMC09wDGDcjtNH7m7KOBj/PkOqykBg4E5Lkkmu2/t4Zn
X5MUkCK4ymm9tHmhWRcBnPEJL/zbGeH9J85rmxYqc5uQ10x9gDxsdxwjY4u8SCsm7GDc82cu7q8T
TAZ14oK+laEGOqmHSn+yoiiHAUuKzYC8Ll/MaOqa+swKAtbMdavXh/aafDQsQk1+4UGrEip7kh5Z
58t2Xje0RsAhGLRunk9x2CaHrD6q754zBVjyEVYFr0pa1yPe7GmcQn+JjuE5D/V/sy+xXbcsjKjy
Klwx322OY2/Cl34LWDMG85LwLP2SWTmwMw8kBIz64xYaSL+WNdhXhaU26fn2qRVkaA2QiulXr4P6
jI5H71jNr25YrZ9qHM/0X++JSMiHJD0cDRDnjtmGIeO3kOR17/JgF5cVB36p66ldFh1ivOuDIJ2l
GMtJJTGniS3QggyNlO5QKrNiWf/OKNWFR0RPWF+f7Gywia43b72OdlvBunZvTE/c6BXjCoq3qAOl
okyW96tz2N8nE/mcEQffQ0LsAhOMpQoq2/zGucNb86AnaUczEx2JVMJorhuX0aIDYpK4r89goKR/
b61iQ0onO51HkzbAn+dcCNwD2yRvndb670bpRbwScfuecoCCAgFfGxhxbmgB0dYaeqRuW2cnDBYZ
APujKaQud51KCO9Jzj2tGuTpQmZSEvvkq3RLJFaTU0Tsj/GevV/Q1qabsLDmR5b5gmYfK/D13SvT
kFStckRtD7iQb/QxquFJEyY5WHhg1BaqMKN5VMvNLcCnBCoHG6ZTiyrOvVSsfcD1R0iv6oDJFVj2
YNBPzUKa/ZTxZXWBS/wfuw9t61+gi5s/QyHdZWvYYj2/FcuPLYaMpEu4AqWT85r5ieB+jWulQudv
Y75eoKdANqtb/OekndV1Kh2nOrvuW92TCI4kK6lH9TC24urfHMgg+1q8LzU2N5LDjrQ4db1ozdoo
RVuPVNyvG+eT5X2J/DmFz8cIFVzLYn6RtmrpSsJRqELGJTnXFT6kRHuQBBjQqGlIaijXBSuYgo5S
deyC1cYjwifxeVlFK8HMp4moZkzApUt192q7JOxC89kHrLl2c/JuKZO3OEyfcS68IZdcngvR6yRP
ofRwu7iWUB5MIEGVZPoMs6eZxXr/bHbyqGfQ+4yck10riRIKp+dm7nnRfTbBnk/in3Ll014OWa7w
o4iZ+2aUI/j3BHgny2Oxta+WM9TY9yBGQ7bsKuRDznxIjmQ3GCfFTpGyqKdsorgx5vI+WPrxNF4Y
nhtTR2HHK5FP+iC+ySipwQtMeZXaVtUj7kn2YhGVsqjLU2GtvBa1SwUiZ9Up9UXfV3oGf6l52HBV
7fCFyOYNWnVDzzPDOjiI7YRYCDJmAQe0Mm7ZDNEGwlvPOOi4SyQOWqT0uh2gSxwSowkSKmjqkKPm
UXdOGbxFDgM2i5o0VDvGDxcab8IaeeBrp3l3IS6LENaZbBzMu3g/fg5RQ6oVc0hLLJfOM4B+fnJf
lBxwSPtpWIclxlVSlbHBY30d2JBc1GRhOJMSGGpTPIeTfJP9piYGqAg/Bq6x/iPXHuoTCcNK2Sb0
GmfhwYEmUL0RUbSkcNa/+xSzIWqk7XKNBDZ+zNYYV2HQvFB20m33eJVCzlCDnAgVLSphyqDToYZE
+xSH+c7jdVhvoWinv4mGpXO/m5UeqkFZsfjV+IchfK54lnLw5QD4RPMXC4HO8tVK6BPeZ0DSUa8g
gAxbf2jtyIKA7cnW3dMEyPFGC9B2trz+zdV68gBQkWoCJDbF5suOYvGC5SGnSga+QHUqu5sVl1DK
upkiHvxI0oDX1VOg1nQR3mjGRPLQsA3PCL1+yM13xL+0cgM17IOgFzXY3qvYXdniYvCR8iKRC9IU
6mXs1HBfBsaI0U6TuMtYR/83NQ8bvdeaoqAOskxzZYEIFEplGt2h8FwE3pAunYJUrb2w7YKEpA9p
bJjkeoWNDa3JV8iS7CoQcfuFlDTKsi3rL9Yta51hK1E27xk2TLQogjbqCboyl4orFWkoItrsoDg/
tr53047kd6E4VWb5V1YW0sTDDo6wY4nZ0L92sfys7fzxm1SeNe9rAFA6xOr01aStbmQX2w68+Nwe
JejfhemsAoC3FThJMVRrHazp9+KDWI6sEeB5c+Dm/QCmO4K5wM8rA8RpypmddSusMYXaO8OJ12np
uepJCHNhF1K67XoMY+HrOEkbCqP2vDWpLAFrcFJ6O71M3Iggw/Uv9nOUtmUfRIpYehZ2LDg5TGKA
E+OffYOvSuX9YskGo2BZBMNMShax4cBktixgY7MWouvdko1jSqxL14+7F0ccVtQhfOcR8mDL4cFJ
E9j6rh1TlVAahTxxS6OPZ3OtcT0XMvV9yciCUgSjMAniYxmnfX5nx77eeqOD1pVMObJASNtD+Jpc
VSUP1Ye9FA08ZIriJJP21yBWbg5/xDlfwDMdkda8wGzEPdP1uxgRgxEqfot4nZc6HBtjPZYXATDY
Dlj6h/hk5CW9G9uXOz3eIGVlC5X/5mWloBgN+rtAXUSYDcHe327SeHJ99khYH6y+ZOt2uJ0by3Fl
yXWWpLN86H+CHs5JZq6poBTS6+GWyuEUW6yh/Uz6gDlwzTuWhuEju+yAw9Px7x7YDcwpfPGFG787
pYeilXv//szbK68qYko/v+cOT2v+0GHq4X/jtDorKriSakc9E3DJdjkgTVbHQbv5Df6Le9fMLPmR
Z6qyPECsu/wvOfaM3beEKxBwTlYvASh7J2vquzuyVA6UwQG64ANtJUVL7VJywkP8wlUdbDKmMBgD
3ev0dhmz2scpG0+T70tycI1Fn9zwQkqRKfVaVHMaqb7xYmIIdsuqlDQq9dHUCnRa1Zb8Hxc6ILCi
LfLsriln6+6OkenP28Zp5xuowZpQBtpThsehokA8felJLFV5uxYG3u617WWSp2/WXZQXj/oUlbzq
j5fIct0pEX7Pzi3iomBMcB3dkSJOPZ4q7mXUABL0Km54m+NWIdBjdCMeejf79eFCeh0BkgsB0OV7
uWHJ4eRuF4iWv27aAQZEZ/jKWxqFVIfO+OlS5hNGV0+72fmF1rVmFYqs9ahWPF4qUZ/qden9lx3H
W8AIXp5elmsO9uuOacc+otAvZR5Luzb0rb2E1dyqWcXFpRVNddv2Nw1BkQnuMMMzHPhC1DCUptsx
hHyRmKPAk+n8nXf7di76YRpVR44F+n8w1wnlvNOTmZi5HhGk1dzKmYShT5yspvYsPzdsv7qw7zv9
DQMjlsUUapQOaTkvNoL0zX9xIzZju4MeIuSfXrwd46wUs3IljL+LLXtfvY9xESJMnu1KTu5/502E
inDhg/RJMxgXNOaatJpBxeGiqFdvzV3IyNYCYOLpzcQCSvRpsHhpkg5mEZAMET6in4Q50RJf/Fvt
oiOsu4fCREIHHXTEKAnQ+lOfNRP0PI4TXym0zzNXWxh8EHfnVOPlJw5krQTmou1Z/Fl7kC1INFzQ
gM1fszwE1xJCPOomAYAO9PX6cJ0hODJYYoEwCMgz1G7QBDgHrYKkT1Fexo83zH/Rcj/cOjXAXWWG
lDUkWRMCr3g7XgY8qiUhiy+pbB8M1rwqZrqobKtiGHjCBkcrBQar2Z8VPO93Fbnx6vEK5vOM/Vsi
56Ppnp8fSdqJGXuYsuJ5sWCDkdwHImD12ahhoAhzsKLBbpHpOh7gkPCgF+f49MuJIBDcpLzrdXT5
HXEqiIu6I0w3cV+x4tPCnpVjvOrqBf+WU2QIRc78ybjy6j3U6sGqSei2yYgCOq55YwM8l0H6uLuF
IAHVpfjIuvtw/sglyu1aTNnwONtMmjQTKWVwQktubBXl9YuJ05KycpJhtNYPilupqJiRreJOyW8o
n6BFm0yPR35rc0BDnKspynO6oS2A+0ihnfr6SXPLOXQCALBbW1TUya1f4/Qvi4I4U1Pym5bHrpY0
Wj6FL8nWnEM87p6l5NhIQkIwvLZ6AxThfGVPXWXnyAI+F3L44LpAPC5f0mtR02uBbTWj4CglrqmQ
d3scaQ2xq8DT0Lv6H3yw5cwupGFYpL5WZpOs/1sFl5TG41x/GPqbkr4FqZx6ui06riZEZxl3JLuY
AbSSqQHiDbguaeH1C9p1xLePxXdU8N1S+TX3lSKyNPMDyVL3QYMisauOChrgUzCjX0AWWB0WIpN9
fEqxSq2ZE/b8BCaOPaU058PN5BKJC8x7kfR5xj0MpyquBFQtGN0M9Fgzp/PP+YzuNSDQOe3TNh5a
o4FT3C/wplW4aOc/WyI0EQXKzeiscYGJIBTXSclQSD+2fWExfcA4a86fpTix7ASy1I86xk0xhyma
WbHyJzVnV8eXtCRhdakprB3BiuepdRpPQgMfn2/3PFiwyLZ1nDDsor72tkjxuJReW//0i1Kqcdpa
Pw9rq/GmLaB45KuRhdLRhHPf9tR83ILbASEXGxQhgi0Y1ZJuuuaGC4xVUud0X1rcQeH11EbCHSqO
amEklFwfJPgCqWRXAF609dsf89XD6rBjcyrUFO+nt0j9LQe2O+hYT5a/pqFjiUta7B0XU9BoQwnL
MKHK8ULDJ9WyDPS6iWvZet/F87ehLC5cY3e5r3thhROJ16CWAGqiNGKpIK96EC7dq8tpdNfJFCGN
1Pgm3QsdxPDMckr2A7O6LgWLQjlM9LVud4QzFnrKcr58WXhFjSNVlPRRMI64WI/SxYnP248wSIIc
kQtLS1XGsBnL7nspRiuSph+VfSZoZk1C2mtnZ5W3xau2TY/dyqQ1jYEk8gIryVsXLHXI0/CCbqA7
vxej/UAT/i3K/nONEADnzG+ono0AvvJQCAlMtbnHj3r0W0clg6huCD3tNr4fzoPb3V9/1CxZ++NV
W3s+fwl7J3htAEuxKawJhyEWhYcK3vXggMEIwi8UWsi4C5Se0vBdND7bIawZ0wWFrNbQaYuJUzYs
AiXKQeLhssZY1eJJLuHqXT7aMBPmSRK8+b+/Cm0b8yIu+FGSnsIzKOybVXJXu3vvtWcLfGyFmSha
ZBExkTTMfWnbcfCCpLhjPXrqIsc+qS5O5GCMkXPP8Kf674KZI38VOPWweCmLztKWHxrT4jS19SFV
jYBkor8l8auP/aWXTL1p4XMFixGcldKgkK9awc02dcH4/XKt0OEnjnGFI9BIOSkNO4eeIH2LpMXR
PwpPMgVfUUcjDtx2CYOExOiqooHiPCAd9URflQgKT2x9FOqkKXfLv1tuX0Xq6JQ50I+kebhGh5zP
8HlxhuWvx4XOYUWH1gWlbdfinrlGwjluttx73qFaMFvZIH8kO6y4k7X6+inX18gfE1lIPKlybCpx
W5tn1swWIYfKQAEqairdxaVAFtt/oURDnoiM1c1HZ5fCn2U1UpK/uXANz2KQJeAVegLf7ojBmE8h
oYVVI3PWVgSQPh9bviX09+/Xu1kx+o6Ax/oR6Yi/WtRm+JLrLQ8qPPJzNmdONsvkh1mvDzs+5gVN
gfIAuyECrJKArkRA+kU+1MJECdNHUkk/pcw00XvK4xVICHHghHNwGQEjISOyUqRDDSOcuCjVWHBt
BNTVVt+nT0mpGmpFMmcOOQN8zkrqr2xMeyZ8KZ0TFro/CMjSqJNZcpsgPqlTvsbkH5ELLyh3U3M3
THIWDOj0HgN04LkxmKVuRBcRH6KibV0Bl+w55KO6HsImBDxSFe3/b2Elc/71gw5C2+7eni5Cryok
GklujTxDjtMHg5pp/Y4alV646OwKcX7us62G8d/6jBSi6cknXQzFlwVOiof5VsWHRFbYzu32skR7
eIgFVei59uunVbrHRFTvLpK/nbDR62nPgWjki+tq1KlDh4t+Ia85RZAYa62Spsu6KwTF4MpfYzQV
QI5U19Kpteft0+PqzXV9kMjt/PDnTrdv+JZh/6bUMJeD8dwf0LpWhyTMw4xO1Y7eVB5gUWSaONkv
9V2vCc/+7OV+i7lVeORQTccNjQ1iibreqkrRzieE4Y30d2YKzx1GfaCGfmBT49j0fbt7Jj/Ije4i
F01vSa8ounlZqgF0tJ1EtfhiL0rw6ZR9gLmNDTRvuCUCkHKU8fBbEnbWVUraDyyHP+GttZSG1BKG
xPc0JRwekIGg+ofst5LWN7UjWNFtl/ebJqp5RulXfNwmGd3kgWRsmE6RAdqkFW5gpn6tGw26ZKJd
McE4SQ4cw9yw62bg8FFvaZEmScG7EE33DW+e+jbyQC5Yc6Of8Us7VCzV8K9GtsLLKF1Y3HM6Y1XJ
+tz0uY9Cm5k3HAPYVlh+CVByoDZJi6M4bsraFibP9yaojmY57Z+ti88CuCt4ggbKKyQyMH8eMK+6
r7OrFlDqBWBFi8Mx5ueLfPg4zOW6DXyoYStWhckmLRqFIb0AaAYhqNYcryo1qO3ryhr6tvSROnZm
ULAQdPR9dDSkPUpLlzY0ReFFH/R6thoKEitAcia6Z1jYPHwKYzozCiXI9ZansSGiKaTryadQcjJo
x8dd4aXoGWiqBTFpB4ImuSGluibMFTOACZa1un4WvkwB/WBf8tEAvdsOrRgQuWgMwou2siluyOpj
NyG5s/QzhdzMbYU/kCDCTWI7JuTjn1A6lg98uD14wexVwjooN9WEolx7308hDK/rYC9PxUj5Vrsd
jo6q05l5mS81YoalO+9GOjR075wu4EIeGZgoKAa8KWr38fQfYZwpjhFXeZybZeVebwX0DC+Xh1St
5TPkLl4Kf3UWiTGcn03oZf1l0g54w3D6SYzigASofPOyjTp+1TFsODKOhD4DL10VEf99J1U9cGHJ
v52iR9siT9KTEx6puS0y1ChYUg47jalhz0H/01VY4iHrk+cBchETHEvkcJvtCLhzDf4J5y1vlzt6
K8LEHqjOTAqip0ybclEJf7/q2/JqfO1RMtCHeOg6v7ghIRZD1OjJPlQBDaNW7By4OVnPY8Pn8CRX
ES2jSE4ujLnUejdPvavnEhzyHWnIRYtM2XkaC5/TzhVcCwaEQmdevVUe1JLwesPW7w97hFAe6WPz
sLbu05ekvq87XaKAj8Q/eKjX6mX4ZjcydSyY2QXTyo26qEa4KUROaJBycoXxZYmNNW2xndPMVtDP
esT50kDHdWQjD+qXQjWfrmL/swilUzbK6JpZIp3J3iAKVdU1ysIaGIRUWDP++Xu3Xv1Ya5/CkCG9
5bwGc6Qtwh5USPRZZdMg3q/dhTl1k79drjDSkLdvxf2xFMEIdj3H0HU6IqBiM2KQircHAcOtRyI0
v1s9zeHtc1AL2aOKsvV7qQOPldfucKKCD3aBv6QIZblizblTQ5Bh1QM0yxDCxtrWJ7zTc0IfJ6EL
tZBFy6wvHu6WAHhxgOssVU7dDrwAdvVIvbec7nY8gEec28N7oGMiKKoLjxk7p2+/dE66RNmFMZmV
gIEKvGh4HAVxgfS/p/o9ALjpXnG6nwnMzBvDehYhnk9PtUjLyl1RKiAUXBvHuZxAfpto7VrFFqsW
w4e+LVfgBd0CNCA1K07TsDjW0P/TYAtROKT0NCgwV2wF6/23BOnYGHwWNu5eWva5tluFT45Rb00r
auXVleK3WMz8jkpfdW2aspjzg95UurFM4F6fweR1FZ9cM+OOz3QcKkut3zUU0ejjLTFf1rMhPxLF
PGYSsQY8rvnJlY0ELPQ6UDR3GEauD0qibBdKkpnU61QuM90LmKOML0cyyIBloV918D2ObU5t+JhN
acke7kQB9qrOppaw7N2s5VqxVkDJWQGxl9RhMI23UR743T/3SBCsJ1uzyaAL3HTh22U/24X/AHt6
n+r4YjZVCkm0FszgmvFooPZu5uMzOTC4UtjHrCKogQwTkVHuejBlFPTt5FAR7GkALide88gvG33j
wro0nZUms5oyLmPIDGr2kqYoV3+vGyAOOVbFG6mmy9RGHdmJR9N6nTcMCPRwGfgRNJqHTuKztpeA
kHtmLhhm0AScec7iAdGbFUwkNTWwiHYSGP1I+r2lDA/P93B85CBbkzFU8oHy+qGDxh0n7HGm7dRr
Oz3cKf7xrxw7taKa3rHrMiZdTBtOLe81mHLathqbNxunQz6BdZM1u8H7g4TbpOpsgYBhHIBsg5KH
v0FsxLkUZNYJ6b533ASLfoqyjHfBdj6NvV46k2nZ2GDs2ieB1GKQtP5S6iBZzEczdo0vfticcsm3
ORbJvyWfxVQaDNy9G1JtNcTd0tEWaNLKTr9IkOOpOF9mwf/ognJq2LqlLogfMmzN5IVVJ8HBPMD2
bTH7hAqVXuPphaoKbwYQHQcx8W+Jmor9c0NHGncpgPQdqVa9w6oLrAjvee3zbX26iyE9NtIGNpwJ
V25xPhNo9OMn5iUww+MY2JdMtDMp4ey6yY1FFXXQ7xyOiN2D1ulwiuwnZj1H1tl6ZV5TjKm8GOlL
+eBPdxW1/qxvz8whMm8FsvaoX7Kazl+0gjW91KgaAY5GzBSPrMoaKy+U8QMv/zrPMxdAsl/khqO1
Ffwcqe0w6MhMTEJYJLa0fQLVkJPcmMAfcVsQi6xWf7n4fQMC/14rXanXUFfV1mCqyoRVKQAQKjwU
2Wce/02nSPUV5vyNPE6yrrku4+gJt2FC3YmvR8RasrhoYMZCPTY4NOXarOYUI78KeIFY1EBj/FIL
ydddrB6dSTAkrcxejodzlzGu5A5f7dgFQ/8//TrH6ZHACsMv7WBIbMcIAH8Ho01o5UQ8obnXsRMy
/4N739SjSjJ6587kDKdCResft5PQcyODbTblVIFP8EQNGKNEsOunWap+uta53hwr066BA+H0Khdn
ekKEUBu8z7eInCsMLfE7sIWhATpXKhEn6M017w/y2o+BPYS0x8qMi8MtYCS+CWIvnuzjVEPP5yDg
q4n03WjebtjZA87J5JPtpCtfgyfYmJtjxUsmXDO9tVefCrJvePiDjbUxlR1waiph6kX1kVb9+FrN
TfNhHmq3WvwgtmvK0BNTqBz58Uz4gsfnAXLkp2jX2DCRvCmNMqgWM17eyq0x+3CQmnYC3+li0Veh
4gwNWLVj7/tSJ6eGdSz+o85Hg86U//6HFCzpizNwQdDGKEd7JcM367qWZjUhpEkrL5lqsG3rt/pL
W4m6GpLuLuxyf48siDxa5uAZ8M9+hT8eN9ks98uTZarjdYX+/6M7rVPYkM0noyeFUx8rUtpdNT2Y
Hus0HWKkLjlxp2ktd64WXoJwo95DKOp5ZygfRMzzBWvQ9/PacDxiTwGOEmTv5AstZzOGSouFYKBO
3yDVUD7fA2Ihg84IGRw/tKxmqPcoyYOZ84ZGcWIjkQtpj8nXQ5XXqky+YqFx4GfXufXev1Cf5zZD
QAh9GqxPVJUcA13MOEDSs5r13yJi0wD81L/I+d0CFAlulZ83tj+CIU+qiqjgfAVX1p/62bILuGjM
px/FB5q/WJ5MenuqFNffEuuMQJRKWJkwIxWe1+YzMVWnG29Ewh8kPORDNlXopGuTrDxXYAHOmPpc
haVsO6Yd10QcaQSRwVINu1YvGtApz5/gnDQYyUkjgu0wwrtTfHk6xmEKcCUmiWtR+Qv6/4Dg0wOW
pcXvD9qk2WVgeFBg+4GAJDf7P+SuRkRDzVewmfrIAXG3xvBQs9tAgBuwn4bvOQ1bTebntgptwCzu
yEmi2X0xyxa5tjPxu9vOdvTlbHSCNWNw9nouNybbOLOIxTlLBmS+uV5lyqOKDM+580BHgEdvCza3
ZeqD+ArpIy/8MwPJ5CTuO8vG0ISmAaVPvvJnznQcTfUYGq825pl84iacBfxmndQ/P/u75tCyxvmu
j1KryUt1Qs8nxpMUqkmHQTPnna5l0HYg2ekc93BRcKPt9Atge3lHE1MKsAY4A9nsFkz+MLJG3wyU
ely1uMONexrTZHBfb6Ln4A/ZCLtdmVNeFIFixyOA2ut2PgMA7KRTdpls4f019XhazqVl1SUBVqxO
R3UH+83AcVK9V9dmOIp1lAIrHdE97oznpNqco/OfnmJEfYbxUNYJIrMm7MmcS15NG8TUoWVQmBsc
U9IQBsH958NcYhCfd1F1zL5HMD2Eo1XC0iZpRxCLzGQP1Uevpi1VNrIGfJGCOunA+DKJmGl1F6wm
uRZ+QDuBZ/TDeN7wgRabC0QhZvH1A6OjZ94nTn9oIqtxZp/9clnhvcgY6Vqr7LHsD27BS6YCFojm
mXKoBnG9Ra7VvvVPbyjw9dFWq3VFAUkBGSFW5Wkoq+34OGwSL8b5idTtFwBqpVd0zEyUqWQzucfI
eH4aVIXq2fit+O7ICJq//Y2bUbZqqmKZgYO3w85Tl/I1cDJoW5ChqicXLABPhhIyIWCMljIA9BD4
oYNh0c/cGf2U7TJvqnidsm9tfeKMvvzQuV90Mmr1PXwmmmbpqS/v9IHwDbM/6e3O98x8NNGzxLXV
YZgg0LOx/fd/khc5P0HmVXHzXrQSxh40xzMz4bwtQRO0V7cqr5kDuugO/0xkhnGz9+6V5AxthSnY
NXSw6Qp0bCAJXT3BuOoShlxMysG3KH9uQMT6FQg0071WHT1g5/4l2K+XrDQQjXVmR8WhaEze9w20
EkMRckAUDXx9TuM453NA3l658NI4zEE3fBDvEUgauckXc2YBfkPH6xHHoOeFLb39b11AqFkwVpMW
PtsFwRpuLOzHMYHRPMP+wSeUI5q/tyfnnWFklRmrAzeaTRQI/lpunI5j3KvnoeCqsu8LPoPcKyLN
+DrKCpWZhss/8OLj6FmgFfCInY9el+XzfzzjD+M9cWCdZbW/Uufsmpmo6OrJ1PTkR5lp7cBjGd62
b4JnxWyaV7vXUsUs+epzaPH0cFRfFc5G5WVVU8RXMXsWM7PfreSBwFhga1koiLBDZnmkZFgv4085
brAvsN7x9xSLgzmjJWs0NZ5OY/w38hGc4GVKuSJSRJpiEIUqeJKtsOYYAQaQuDsqJmSYXiSpBgtM
6FU/D+jd+l23SDW4BRQkJ2WstoHC1SXHZ8Br4MujJ1TCWqPmwW4AsCQeb/7UESuYUH1OTI70TfxJ
nylCZdlPclO2mx4I5hsJvH/UdbRP9uCTTOzmgBlkQXq7nm5JOEyqUhl48KVEDcCPXTY93Gr60Kfo
4qzBmb9VWuZtSEZ3D7MmcpJjjnTihMyD+CDJgB22GZGcllKYkEfN8JzhrUS8w1QQg5+iklB0W8q0
ljnmS70c5qfBVPitETtG7xlia++yP55CrEhsg5VAVR/vGoKKaFxPmME0+ZwNf1053Z7fBEvxl4IU
9TRfWVcTvl8eluGNCHJuhR0bDV4giV+AiUB0oz270Jgg4BobX74Zoa15Dskx26jYYvrQTZPOThbb
7kUgmhURTylE14tVzYlPi2Ion6PDpmKICv3tDthM6OahJmV60UZSI/F3UIWJp1VZmL9WfSUJ5Sv2
oCJbcQgVwFCqKbfI36RfG5+bQGEe35gTPKe3b63odIXBqjSSodX9GFv99paiR+/L1f9ESuisDPTu
EPOoAMRfx+CzDAFOnfuylwt2Jd5/Kt+4C24frcKVRtSA69jBpCV3/r8bO85JSe8xlLrstvr0MvZP
9Zqz5iAb/Dx1+sFtcq/jFLrga+V3P/WukqEAe23/KCxaj20sCLsthLTafTP6dhc7J/VnmjsVqP2R
91W8wagYVO4OfBmW0JSH/NJnEYGWr7YO9icddaIOSCP0HP21QXJtlLrWI9TSalyuuySnEh/oVBQC
gp7MyoV3LCDyLrUkjulrhiNlrTenxR8XxK0Berfh9AKZPzBtEl/eZoHbHhyC4IppTBolF//JNtkN
qLMjdj4YHY2xPjLGY32piSjTzHnv5yz5iYdDLhFL+QnTvixspFkVg/9BUB+L4qaBOo9TUYJ/pTRx
7D06cxvG4ZuzaYS/SBDresWyFg1/EXIoKdfGeH72xMgDncsrtwv5/QyHwmldQ6b+LnsEcKezuf+x
YtC7DxIzOXzhtTCrYQ/OinkWMxrUPysaLoX7BRISy0e+WnpN+6B1Si41Wgr3dEHwPn2ILvlbs5Vp
RjX8gw81HvP7eI3iubMdB5HKOvsfc/fqPCwzmGf8VdacP9chtR1l8olZN3Ue/FHKIFEZnri9LVBL
oEaA0OwBgru9wLQqrZP4HfDsHaUO2/r/gXaaXb96ql3YLDxTE9wRg/TrRDGof53NM/mf0l8+pCUu
3a5NR+Bji7SkRGuxMpx5KKAWPSPsGRjk6uusWZKgGJQN5Ej5+Cw6uVPIxTjSDh2ocLLO2EgPH7F8
bofPQ+Ge/g4gk0lDXMsrEM6iUbM/juGWkgBjOmbhHuJyu0Hbctr9QkaUHVtLQs4uLKlP/c7DnKMD
Vut0fZR8BL/z6x5EHCd2kLN2USadGGli57b1BmImSRvvjo+bpJIKMADwYFb6kismpVG2pwFlBj8E
FSBb8Bz/73vrYe8ynuDU0gYsn9tt3RecRuHkFipzQdG1PZoO6gQgKoD9v/Gq8lnGcBSZxzGWAhse
YizBBE9fqMsFiA6ue00nh1CiByySYR02tsSmnCp6kPuL+4UhmG1U4a9OaC368yshPaGAkK5l9iXz
B5f4d05KbIFGI01fMlHACaldAc+uXVQfYElvYuKu+M0M9I0C1qvmuk8wEW6Q4uM8KxfNV8QwATVk
OfSkz69RZb4Yrqc0AzGqJ15N7Dq8WyHd6oR92FOC3+d4n14wMVXNHvdry5s/5R60Hi/3IyjuPAdf
a0RwqXwNgWDAi+GAOZZht1orA9OfZFkoiyYwYXgMICFGbdpsbdiX/FrxIVnf55EJQC3rnmqTL3lV
otcRWZQygWNiPz8chkMhwvfUeXIjwgyBiUJcs3rZf7H8d4E5nyv0aIRjbCkaGPE9yUdb19rspARJ
gXj6qPcbRDeXmdMz4aZIHuH+KqdeyXB5bC3KjSyQe23KqQBf71406TTkewW64eEDbmGvwxU6G8lZ
/0NgK3W5+wyY45kPgkgrJZ4NkGZL551G2wzO/KBRpa4sl4HKulSKWA0OSCuafPREsv3UFPikQBUB
k7TNp1IQ+C5gXDCDNPV8gUCiljnUfjdbxLO9MGvBOFDmhTJf/jDwCAJD3UNHRFiSNBP4bqajWCTc
O3wr9gS8prF1Ql9yf+RWjrVWRoggozUADwtNfZMpdEZFKJKGwhTFO5rKUgQnvyyWjmSTIoEt0I0r
jlUch8TRXXo+I0Nmc5gC7nqvlNbz+1P7HjxUqAne8zLmggAJ/acnLam6pggMaDHbdAK61O1l7Xk6
T5v1cO0F+FMtuScnPRHvGdVgyS5DXDBWoN6/R38wkapGf/iAOZZryQV3Khog+eqgcYHLvmW4n2vn
9nuf7FCl+Wzf0/WYBvCBYzTH6v66j4Saw29Gy4UuA8Blsl0IHO4NpQsZz52tDvtxEIRC9/wsAy2g
8XKBMQ+FdEClEh8sLX2FepHv3ywdyKaSNW+8vKeOzJELRWCaPhBmyjcJguUtfBRAVq5NfMEMQ+rR
r+wN30wuGQfijNmmyPdMRPARjkT+auPErsb35+B36y1NpHvuRqMHihkwVtV4g/zDfZwLRYfn8ThA
cURBfI4vHAu4oFgsmnYtnUpJW3LkSAOjE8MXfkGE5EC84KaDJMoNW6XS8zEuo8WJIqo00rOlPiNL
93rMsG7u4b9Oh+QMA+4trDLNZedxElYMt5a/x311YPAzlPHhduVAtwMWYPRY52j38nHdWAWVbbf7
g6JENXsIxiM/RtS9osKwJQBavz0ej2R3bGtYULJEiEAecgc+0auoh5ixQxh5a05G9R0IpuC8hP3T
Z6FB9ZiHtCiLb9GWmosFASI/wy5gr0WtRWkHFlh6ZAq4qiytqt8uCeMOvZRgHn3F4y7k809QZdqG
0zYMTO71erOG1tVzBj4xy34j+dX9mhZuxDsAvSqK3YTJ/3Bd6NvGR47NQCrwBwK9lrwI4+HWWoiK
eUnPcawK7pvE06eezncmgQ8z3Zd15Y+557fS2nMgqH9ILL3OUNWmEBfw7LJqB09nsKMdWCvPBaZl
zxslhrV2qkFukKKdrSvQSQMV2ySb1c5XFSwKWtyInh1u9fVu7ArdShFCE5wjM0byO9snqj4dwRxc
bD0hCAA14arOVxWUHB8CiCDnaa/mTEf7J8RK9QF/n52H9wzYQLCcDZXMk8lFQaE3YXUNJ1Xyw6mJ
zn47cgZpDoQBD4iGfDQHdLOq3gF+J6s1oFkqOyehr2siRdaOyUBfF64bz7zKx2Q5L+w2uQBNe48u
6ScT1AT/up4KIejqGUZuSbbAVEzi+e5AeF/0VxaAUxlheyZCcytWRK0xntLojglu3dxqF8aCaA2R
Yto94Fjoo8feGy3Qz21JxtejJTsGgILZL16ybD6tWCM1uW79T4fuYo45M5xHw8O2xqvYCECUh0t4
UJMZ0HNUWOuPbT5Mef7pS3wmkSP3Uxl1K6SCe4gPvrBLgctdKbHShZDAucX245Rmvm5xnrgKJv+8
wHNOBvBjLzQM2vkYNmnUNDfSE4taWQrNChUNbMSG3MTU75rzTmmtAlZuQN0Vv2yLD2yGd2rqSdt+
ArrGTVzEBFF4OuYpQ6hVdHSoRIHDFrFLXkHCad49Q7bsibPOQmU865cKYWU9b0Ba+K5hBo7+yXcZ
qR6ZWrGoyvkbX9tLelvT0msFcXxbPdYVvHsCBVsJ400X92v+gYJFPJKaMjFtoJjB7to403nl3df4
poQDh39te4W62h5JadSPBEU3YqP7IWBNLYUvRE835WA+rBpysxXVAui5IC5f22wcdfdelr80iOkS
`protect end_protected
