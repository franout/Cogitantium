module compact_and_select ();

endmodule