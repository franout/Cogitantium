// Register NVDLA_SDP_S_STATUS_0
#define NVDLA_SDP_S_STATUS_0					32'h9000
#define NVDLA_SDP_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_SDP_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_SDP_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_SDP_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_SDP_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_SDP_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_SDP_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_SDP_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_SDP_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_SDP_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_SDP_S_POINTER_0
#define NVDLA_SDP_S_POINTER_0					32'h9004
#define NVDLA_SDP_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_SDP_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_SDP_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_SDP_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_SDP_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_SDP_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_SDP_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_SDP_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_SDP_S_LUT_ACCESS_CFG_0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0					32'h9008
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ADDR_RANGE			9:0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ADDR_SIZE				10
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_RANGE			16:16
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_SIZE				1
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_LE			1'h0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_TABLE_ID_LO			1'h1
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_RANGE			17:17
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_SIZE				1
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_READ			1'h0
#define NVDLA_SDP_S_LUT_ACCESS_CFG_0_LUT_ACCESS_TYPE_WRITE			1'h1


// Register NVDLA_SDP_S_LUT_ACCESS_DATA_0
#define NVDLA_SDP_S_LUT_ACCESS_DATA_0					32'h900c
#define NVDLA_SDP_S_LUT_ACCESS_DATA_0_LUT_DATA_RANGE			15:0
#define NVDLA_SDP_S_LUT_ACCESS_DATA_0_LUT_DATA_SIZE				16


// Register NVDLA_SDP_S_LUT_CFG_0
#define NVDLA_SDP_S_LUT_CFG_0					32'h9010
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_RANGE			0:0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_EXPONENT			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_LE_FUNCTION_LINEAR			1'h1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_RANGE			4:4
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_LE			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_UFLOW_PRIORITY_LO			1'h1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_RANGE			5:5
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_LE			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_OFLOW_PRIORITY_LO			1'h1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_RANGE			6:6
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_SIZE				1
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_LE			1'h0
#define NVDLA_SDP_S_LUT_CFG_0_LUT_HYBRID_PRIORITY_LO			1'h1


// Register NVDLA_SDP_S_LUT_INFO_0
#define NVDLA_SDP_S_LUT_INFO_0					32'h9014
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_OFFSET_RANGE			7:0
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_OFFSET_SIZE				8
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_SELECT_RANGE			15:8
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LE_INDEX_SELECT_SIZE				8
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LO_INDEX_SELECT_RANGE			23:16
#define NVDLA_SDP_S_LUT_INFO_0_LUT_LO_INDEX_SELECT_SIZE				8


// Register NVDLA_SDP_S_LUT_LE_START_0
#define NVDLA_SDP_S_LUT_LE_START_0					32'h9018
#define NVDLA_SDP_S_LUT_LE_START_0_LUT_LE_START_RANGE			31:0
#define NVDLA_SDP_S_LUT_LE_START_0_LUT_LE_START_SIZE				32


// Register NVDLA_SDP_S_LUT_LE_END_0
#define NVDLA_SDP_S_LUT_LE_END_0					32'h901c
#define NVDLA_SDP_S_LUT_LE_END_0_LUT_LE_END_RANGE			31:0
#define NVDLA_SDP_S_LUT_LE_END_0_LUT_LE_END_SIZE				32


// Register NVDLA_SDP_S_LUT_LO_START_0
#define NVDLA_SDP_S_LUT_LO_START_0					32'h9020
#define NVDLA_SDP_S_LUT_LO_START_0_LUT_LO_START_RANGE			31:0
#define NVDLA_SDP_S_LUT_LO_START_0_LUT_LO_START_SIZE				32


// Register NVDLA_SDP_S_LUT_LO_END_0
#define NVDLA_SDP_S_LUT_LO_END_0					32'h9024
#define NVDLA_SDP_S_LUT_LO_END_0_LUT_LO_END_RANGE			31:0
#define NVDLA_SDP_S_LUT_LO_END_0_LUT_LO_END_SIZE				32


// Register NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0					32'h9028
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_UFLOW_SCALE_RANGE			15:0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_UFLOW_SCALE_SIZE				16
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_OFLOW_SCALE_RANGE			31:16
#define NVDLA_SDP_S_LUT_LE_SLOPE_SCALE_0_LUT_LE_SLOPE_OFLOW_SCALE_SIZE				16


// Register NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0					32'h902c
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_UFLOW_SHIFT_RANGE			4:0
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_UFLOW_SHIFT_SIZE				5
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_OFLOW_SHIFT_RANGE			9:5
#define NVDLA_SDP_S_LUT_LE_SLOPE_SHIFT_0_LUT_LE_SLOPE_OFLOW_SHIFT_SIZE				5


// Register NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0					32'h9030
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_UFLOW_SCALE_RANGE			15:0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_UFLOW_SCALE_SIZE				16
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_OFLOW_SCALE_RANGE			31:16
#define NVDLA_SDP_S_LUT_LO_SLOPE_SCALE_0_LUT_LO_SLOPE_OFLOW_SCALE_SIZE				16


// Register NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0					32'h9034
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_UFLOW_SHIFT_RANGE			4:0
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_UFLOW_SHIFT_SIZE				5
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_OFLOW_SHIFT_RANGE			9:5
#define NVDLA_SDP_S_LUT_LO_SLOPE_SHIFT_0_LUT_LO_SLOPE_OFLOW_SHIFT_SIZE				5


// Register NVDLA_SDP_D_OP_ENABLE_0
#define NVDLA_SDP_D_OP_ENABLE_0					32'h9038
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_SDP_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_SDP_D_DATA_CUBE_WIDTH_0
#define NVDLA_SDP_D_DATA_CUBE_WIDTH_0					32'h903c
#define NVDLA_SDP_D_DATA_CUBE_WIDTH_0_WIDTH_RANGE			12:0
#define NVDLA_SDP_D_DATA_CUBE_WIDTH_0_WIDTH_SIZE				13


// Register NVDLA_SDP_D_DATA_CUBE_HEIGHT_0
#define NVDLA_SDP_D_DATA_CUBE_HEIGHT_0					32'h9040
#define NVDLA_SDP_D_DATA_CUBE_HEIGHT_0_HEIGHT_RANGE			12:0
#define NVDLA_SDP_D_DATA_CUBE_HEIGHT_0_HEIGHT_SIZE				13


// Register NVDLA_SDP_D_DATA_CUBE_CHANNEL_0
#define NVDLA_SDP_D_DATA_CUBE_CHANNEL_0					32'h9044
#define NVDLA_SDP_D_DATA_CUBE_CHANNEL_0_CHANNEL_RANGE			12:0
#define NVDLA_SDP_D_DATA_CUBE_CHANNEL_0_CHANNEL_SIZE				13


// Register NVDLA_SDP_D_DST_BASE_ADDR_LOW_0
#define NVDLA_SDP_D_DST_BASE_ADDR_LOW_0					32'h9048
#define NVDLA_SDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_SDP_D_DST_BASE_ADDR_LOW_0_DST_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0
#define NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0					32'h904c
#define NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_SDP_D_DST_BASE_ADDR_HIGH_0_DST_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_SDP_D_DST_LINE_STRIDE_0
#define NVDLA_SDP_D_DST_LINE_STRIDE_0					32'h9050
#define NVDLA_SDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_RANGE			31:0
#define NVDLA_SDP_D_DST_LINE_STRIDE_0_DST_LINE_STRIDE_SIZE				32


// Register NVDLA_SDP_D_DST_SURFACE_STRIDE_0
#define NVDLA_SDP_D_DST_SURFACE_STRIDE_0					32'h9054
#define NVDLA_SDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_SDP_D_DST_SURFACE_STRIDE_0_DST_SURFACE_STRIDE_SIZE				32


// Register NVDLA_SDP_D_DP_BS_CFG_0
#define NVDLA_SDP_D_DP_BS_CFG_0					32'h9058
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_RANGE			0:0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_RANGE			3:2
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_SIZE				2
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_MAX			2'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_MIN			2'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_ALU_ALGO_SUM			2'h2
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_RANGE			4:4
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_RANGE			5:5
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_MUL_PRELU_YES			1'h1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_RANGE			6:6
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BS_CFG_0_BS_RELU_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_BS_ALU_CFG_0
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0					32'h905c
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SHIFT_VALUE_RANGE			13:8
#define NVDLA_SDP_D_DP_BS_ALU_CFG_0_BS_ALU_SHIFT_VALUE_SIZE				6


// Register NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0					32'h9060
#define NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0_BS_ALU_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BS_ALU_SRC_VALUE_0_BS_ALU_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_BS_MUL_CFG_0
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0					32'h9064
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SHIFT_VALUE_RANGE			15:8
#define NVDLA_SDP_D_DP_BS_MUL_CFG_0_BS_MUL_SHIFT_VALUE_SIZE				8


// Register NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0					32'h9068
#define NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0_BS_MUL_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BS_MUL_SRC_VALUE_0_BS_MUL_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_BN_CFG_0
#define NVDLA_SDP_D_DP_BN_CFG_0					32'h906c
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_RANGE			0:0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_RANGE			3:2
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_SIZE				2
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_MAX			2'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_MIN			2'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_ALU_ALGO_SUM			2'h2
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_RANGE			4:4
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_RANGE			5:5
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_MUL_PRELU_YES			1'h1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_RANGE			6:6
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_BN_CFG_0_BN_RELU_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_BN_ALU_CFG_0
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0					32'h9070
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SHIFT_VALUE_RANGE			13:8
#define NVDLA_SDP_D_DP_BN_ALU_CFG_0_BN_ALU_SHIFT_VALUE_SIZE				6


// Register NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0					32'h9074
#define NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0_BN_ALU_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BN_ALU_SRC_VALUE_0_BN_ALU_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_BN_MUL_CFG_0
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0					32'h9078
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_SIZE				1
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SHIFT_VALUE_RANGE			15:8
#define NVDLA_SDP_D_DP_BN_MUL_CFG_0_BN_MUL_SHIFT_VALUE_SIZE				8


// Register NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0
#define NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0					32'h907c
#define NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0_BN_MUL_OPERAND_RANGE			15:0
#define NVDLA_SDP_D_DP_BN_MUL_SRC_VALUE_0_BN_MUL_OPERAND_SIZE				16


// Register NVDLA_SDP_D_DP_EW_CFG_0
#define NVDLA_SDP_D_DP_EW_CFG_0					32'h9080
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_RANGE			0:0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_RANGE			3:2
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_SIZE				2
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_MAX			2'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_MIN			2'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_SUM			2'h2
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_ALU_ALGO_EQL			2'h3
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_RANGE			4:4
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_BYPASS_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_RANGE			5:5
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_MUL_PRELU_YES			1'h1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_RANGE			6:6
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_CFG_0_EW_LUT_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_EW_ALU_CFG_0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0					32'h9084
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_SIZE				1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_ALU_CFG_0_EW_ALU_CVT_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0					32'h9088
#define NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0_EW_ALU_OPERAND_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_ALU_SRC_VALUE_0_EW_ALU_OPERAND_SIZE				32


// Register NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0					32'h908c
#define NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0_EW_ALU_CVT_OFFSET_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_OFFSET_VALUE_0_EW_ALU_CVT_OFFSET_SIZE				32


// Register NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0					32'h9090
#define NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0_EW_ALU_CVT_SCALE_RANGE			15:0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_SCALE_VALUE_0_EW_ALU_CVT_SCALE_SIZE				16


// Register NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0					32'h9094
#define NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0_EW_ALU_CVT_TRUNCATE_RANGE			5:0
#define NVDLA_SDP_D_DP_EW_ALU_CVT_TRUNCATE_VALUE_0_EW_ALU_CVT_TRUNCATE_SIZE				6


// Register NVDLA_SDP_D_DP_EW_MUL_CFG_0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0					32'h9098
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_RANGE			0:0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_SIZE				1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_REG			1'h0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_SRC_MEM			1'h1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_RANGE			1:1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_SIZE				1
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_NO			1'h0
#define NVDLA_SDP_D_DP_EW_MUL_CFG_0_EW_MUL_CVT_BYPASS_YES			1'h1


// Register NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0					32'h909c
#define NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0_EW_MUL_OPERAND_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_MUL_SRC_VALUE_0_EW_MUL_OPERAND_SIZE				32


// Register NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0					32'h90a0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0_EW_MUL_CVT_OFFSET_RANGE			31:0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_OFFSET_VALUE_0_EW_MUL_CVT_OFFSET_SIZE				32


// Register NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0					32'h90a4
#define NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0_EW_MUL_CVT_SCALE_RANGE			15:0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_SCALE_VALUE_0_EW_MUL_CVT_SCALE_SIZE				16


// Register NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0					32'h90a8
#define NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0_EW_MUL_CVT_TRUNCATE_RANGE			5:0
#define NVDLA_SDP_D_DP_EW_MUL_CVT_TRUNCATE_VALUE_0_EW_MUL_CVT_TRUNCATE_SIZE				6


// Register NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0
#define NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0					32'h90ac
#define NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0_EW_TRUNCATE_RANGE			9:0
#define NVDLA_SDP_D_DP_EW_TRUNCATE_VALUE_0_EW_TRUNCATE_SIZE				10


// Register NVDLA_SDP_D_FEATURE_MODE_CFG_0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0					32'h90b0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_RANGE			0:0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_OFF			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_FLYING_MODE_ON			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_RANGE			1:1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_MEM			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_OUTPUT_DST_PDP			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_RANGE			2:2
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_OFF			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_WINOGRAD_ON			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_RANGE			3:3
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_SIZE				1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_DISABLE			1'h0
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_NAN_TO_ZERO_ENABLE			1'h1
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_RANGE			12:8
#define NVDLA_SDP_D_FEATURE_MODE_CFG_0_BATCH_NUMBER_SIZE				5


// Register NVDLA_SDP_D_DST_DMA_CFG_0
#define NVDLA_SDP_D_DST_DMA_CFG_0					32'h90b4
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_RANGE			0:0
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_SIZE				1
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_CV			1'h0
#define NVDLA_SDP_D_DST_DMA_CFG_0_DST_RAM_TYPE_MC			1'h1


// Register NVDLA_SDP_D_DST_BATCH_STRIDE_0
#define NVDLA_SDP_D_DST_BATCH_STRIDE_0					32'h90b8
#define NVDLA_SDP_D_DST_BATCH_STRIDE_0_DST_BATCH_STRIDE_RANGE			31:0
#define NVDLA_SDP_D_DST_BATCH_STRIDE_0_DST_BATCH_STRIDE_SIZE				32


// Register NVDLA_SDP_D_DATA_FORMAT_0
#define NVDLA_SDP_D_DATA_FORMAT_0					32'h90bc
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_RANGE			1:0
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_SIZE				2
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_SDP_D_DATA_FORMAT_0_PROC_PRECISION_FP16			2'h2
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_RANGE			3:2
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_SIZE				2
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_INT8			2'h0
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_INT16			2'h1
#define NVDLA_SDP_D_DATA_FORMAT_0_OUT_PRECISION_FP16			2'h2


// Register NVDLA_SDP_D_CVT_OFFSET_0
#define NVDLA_SDP_D_CVT_OFFSET_0					32'h90c0
#define NVDLA_SDP_D_CVT_OFFSET_0_CVT_OFFSET_RANGE			31:0
#define NVDLA_SDP_D_CVT_OFFSET_0_CVT_OFFSET_SIZE				32


// Register NVDLA_SDP_D_CVT_SCALE_0
#define NVDLA_SDP_D_CVT_SCALE_0					32'h90c4
#define NVDLA_SDP_D_CVT_SCALE_0_CVT_SCALE_RANGE			15:0
#define NVDLA_SDP_D_CVT_SCALE_0_CVT_SCALE_SIZE				16


// Register NVDLA_SDP_D_CVT_SHIFT_0
#define NVDLA_SDP_D_CVT_SHIFT_0					32'h90c8
#define NVDLA_SDP_D_CVT_SHIFT_0_CVT_SHIFT_RANGE			5:0
#define NVDLA_SDP_D_CVT_SHIFT_0_CVT_SHIFT_SIZE				6


// Register NVDLA_SDP_D_STATUS_0
#define NVDLA_SDP_D_STATUS_0					32'h90cc
#define NVDLA_SDP_D_STATUS_0_STATUS_UNEQUAL_RANGE			0:0
#define NVDLA_SDP_D_STATUS_0_STATUS_UNEQUAL_SIZE				1


// Register NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0
#define NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0					32'h90d0
#define NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_D_STATUS_NAN_INPUT_NUM_0_STATUS_NAN_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0
#define NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0					32'h90d4
#define NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_RANGE			31:0
#define NVDLA_SDP_D_STATUS_INF_INPUT_NUM_0_STATUS_INF_INPUT_NUM_SIZE				32


// Register NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0
#define NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0					32'h90d8
#define NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0_STATUS_NAN_OUTPUT_NUM_RANGE			31:0
#define NVDLA_SDP_D_STATUS_NAN_OUTPUT_NUM_0_STATUS_NAN_OUTPUT_NUM_SIZE				32


// Register NVDLA_SDP_D_PERF_ENABLE_0
#define NVDLA_SDP_D_PERF_ENABLE_0					32'h90dc
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_RANGE			0:0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_DMA_EN_YES			1'h1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_RANGE			1:1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_LUT_EN_YES			1'h1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_RANGE			2:2
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_SAT_EN_YES			1'h1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_RANGE			3:3
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_SIZE				1
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_NO			1'h0
#define NVDLA_SDP_D_PERF_ENABLE_0_PERF_NAN_INF_COUNT_EN_YES			1'h1


// Register NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0
#define NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0					32'h90e0
#define NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0_WDMA_STALL_RANGE			31:0
#define NVDLA_SDP_D_PERF_WDMA_WRITE_STALL_0_WDMA_STALL_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_UFLOW_0
#define NVDLA_SDP_D_PERF_LUT_UFLOW_0					32'h90e4
#define NVDLA_SDP_D_PERF_LUT_UFLOW_0_LUT_UFLOW_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_UFLOW_0_LUT_UFLOW_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_OFLOW_0
#define NVDLA_SDP_D_PERF_LUT_OFLOW_0					32'h90e8
#define NVDLA_SDP_D_PERF_LUT_OFLOW_0_LUT_OFLOW_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_OFLOW_0_LUT_OFLOW_SIZE				32


// Register NVDLA_SDP_D_PERF_OUT_SATURATION_0
#define NVDLA_SDP_D_PERF_OUT_SATURATION_0					32'h90ec
#define NVDLA_SDP_D_PERF_OUT_SATURATION_0_OUT_SATURATION_RANGE			31:0
#define NVDLA_SDP_D_PERF_OUT_SATURATION_0_OUT_SATURATION_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_HYBRID_0
#define NVDLA_SDP_D_PERF_LUT_HYBRID_0					32'h90f0
#define NVDLA_SDP_D_PERF_LUT_HYBRID_0_LUT_HYBRID_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_HYBRID_0_LUT_HYBRID_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_LE_HIT_0
#define NVDLA_SDP_D_PERF_LUT_LE_HIT_0					32'h90f4
#define NVDLA_SDP_D_PERF_LUT_LE_HIT_0_LUT_LE_HIT_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_LE_HIT_0_LUT_LE_HIT_SIZE				32


// Register NVDLA_SDP_D_PERF_LUT_LO_HIT_0
#define NVDLA_SDP_D_PERF_LUT_LO_HIT_0					32'h90f8
#define NVDLA_SDP_D_PERF_LUT_LO_HIT_0_LUT_LO_HIT_RANGE			31:0
#define NVDLA_SDP_D_PERF_LUT_LO_HIT_0_LUT_LO_HIT_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_SDP	32'h9000
