// Register NVDLA_GLB_S_NVDLA_HW_VERSION_0
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0					32'h1000
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MAJOR_RANGE			7:0
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MAJOR_SIZE				8
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MINOR_RANGE			23:8
#define NVDLA_GLB_S_NVDLA_HW_VERSION_0_MINOR_SIZE				16


// Register NVDLA_GLB_S_INTR_MASK_0
#define NVDLA_GLB_S_INTR_MASK_0					32'h1004
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK0_RANGE			0:0
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK1_RANGE			1:1
#define NVDLA_GLB_S_INTR_MASK_0_SDP_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK0_RANGE			2:2
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK1_RANGE			3:3
#define NVDLA_GLB_S_INTR_MASK_0_CDP_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK0_RANGE			4:4
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK1_RANGE			5:5
#define NVDLA_GLB_S_INTR_MASK_0_PDP_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK0_RANGE			6:6
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK1_RANGE			7:7
#define NVDLA_GLB_S_INTR_MASK_0_BDMA_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK0_RANGE			8:8
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK1_RANGE			9:9
#define NVDLA_GLB_S_INTR_MASK_0_RUBIK_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK0_RANGE			16:16
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK1_RANGE			17:17
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_DAT_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK0_RANGE			18:18
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK1_RANGE			19:19
#define NVDLA_GLB_S_INTR_MASK_0_CDMA_WT_DONE_MASK1_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK0_RANGE			20:20
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK0_SIZE				1
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK1_RANGE			21:21
#define NVDLA_GLB_S_INTR_MASK_0_CACC_DONE_MASK1_SIZE				1


// Register NVDLA_GLB_S_INTR_SET_0
#define NVDLA_GLB_S_INTR_SET_0					32'h1008
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET0_RANGE			0:0
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET1_RANGE			1:1
#define NVDLA_GLB_S_INTR_SET_0_SDP_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET0_RANGE			2:2
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET1_RANGE			3:3
#define NVDLA_GLB_S_INTR_SET_0_CDP_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET0_RANGE			4:4
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET1_RANGE			5:5
#define NVDLA_GLB_S_INTR_SET_0_PDP_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET0_RANGE			6:6
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET1_RANGE			7:7
#define NVDLA_GLB_S_INTR_SET_0_BDMA_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET0_RANGE			8:8
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET1_RANGE			9:9
#define NVDLA_GLB_S_INTR_SET_0_RUBIK_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET0_RANGE			16:16
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET1_RANGE			17:17
#define NVDLA_GLB_S_INTR_SET_0_CDMA_DAT_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET0_RANGE			18:18
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET1_RANGE			19:19
#define NVDLA_GLB_S_INTR_SET_0_CDMA_WT_DONE_SET1_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET0_RANGE			20:20
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET0_SIZE				1
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET1_RANGE			21:21
#define NVDLA_GLB_S_INTR_SET_0_CACC_DONE_SET1_SIZE				1


// Register NVDLA_GLB_S_INTR_STATUS_0
#define NVDLA_GLB_S_INTR_STATUS_0					32'h100c
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS0_RANGE			0:0
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS1_RANGE			1:1
#define NVDLA_GLB_S_INTR_STATUS_0_SDP_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS0_RANGE			2:2
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS1_RANGE			3:3
#define NVDLA_GLB_S_INTR_STATUS_0_CDP_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS0_RANGE			4:4
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS1_RANGE			5:5
#define NVDLA_GLB_S_INTR_STATUS_0_PDP_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS0_RANGE			6:6
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS1_RANGE			7:7
#define NVDLA_GLB_S_INTR_STATUS_0_BDMA_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS0_RANGE			8:8
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS1_RANGE			9:9
#define NVDLA_GLB_S_INTR_STATUS_0_RUBIK_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS0_RANGE			16:16
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS1_RANGE			17:17
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_DAT_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS0_RANGE			18:18
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS1_RANGE			19:19
#define NVDLA_GLB_S_INTR_STATUS_0_CDMA_WT_DONE_STATUS1_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS0_RANGE			20:20
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS0_SIZE				1
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS1_RANGE			21:21
#define NVDLA_GLB_S_INTR_STATUS_0_CACC_DONE_STATUS1_SIZE				1



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_GLB	32'h1000
