// Register NVDLA_PDP_RDMA_S_STATUS_0
#define NVDLA_PDP_RDMA_S_STATUS_0					32'ha000
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_PDP_RDMA_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_PDP_RDMA_S_POINTER_0
#define NVDLA_PDP_RDMA_S_POINTER_0					32'ha004
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_PDP_RDMA_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_PDP_RDMA_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_PDP_RDMA_D_OP_ENABLE_0
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0					32'ha008
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_PDP_RDMA_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0					32'ha00c
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_RANGE			12:0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_WIDTH_0_CUBE_IN_WIDTH_SIZE				13


// Register NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0					32'ha010
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_RANGE			12:0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_HEIGHT_0_CUBE_IN_HEIGHT_SIZE				13


// Register NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0					32'ha014
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_RANGE			12:0
#define NVDLA_PDP_RDMA_D_DATA_CUBE_IN_CHANNEL_0_CUBE_IN_CHANNEL_SIZE				13


// Register NVDLA_PDP_RDMA_D_FLYING_MODE_0
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0					32'ha018
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_RANGE			0:0
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_SIZE				1
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_ON_FLYING			1'h0
#define NVDLA_PDP_RDMA_D_FLYING_MODE_0_FLYING_MODE_OFF_FLYING			1'h1


// Register NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0					32'ha01c
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_LOW_0_SRC_BASE_ADDR_LOW_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0					32'ha020
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_BASE_ADDR_HIGH_0_SRC_BASE_ADDR_HIGH_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0
#define NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0					32'ha024
#define NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_LINE_STRIDE_0_SRC_LINE_STRIDE_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0
#define NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0					32'ha028
#define NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_RANGE			31:0
#define NVDLA_PDP_RDMA_D_SRC_SURFACE_STRIDE_0_SRC_SURFACE_STRIDE_SIZE				32


// Register NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0					32'ha02c
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_RANGE			0:0
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_SIZE				1
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_CV			1'h0
#define NVDLA_PDP_RDMA_D_SRC_RAM_CFG_0_SRC_RAM_TYPE_MC			1'h1


// Register NVDLA_PDP_RDMA_D_DATA_FORMAT_0
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0					32'ha030
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_RANGE			1:0
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_SIZE				2
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_INT8			2'h0
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_INT16			2'h1
#define NVDLA_PDP_RDMA_D_DATA_FORMAT_0_INPUT_DATA_FP16			2'h2


// Register NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0
#define NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0					32'ha034
#define NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0_SPLIT_NUM_RANGE			7:0
#define NVDLA_PDP_RDMA_D_OPERATION_MODE_CFG_0_SPLIT_NUM_SIZE				8


// Register NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0					32'ha038
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_RANGE			3:0
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_SIZE				4
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_1			4'h0
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_2			4'h1
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_3			4'h2
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_4			4'h3
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_5			4'h4
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_6			4'h5
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_7			4'h6
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_WIDTH_KERNEL_WIDTH_8			4'h7
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_RANGE			7:4
#define NVDLA_PDP_RDMA_D_POOLING_KERNEL_CFG_0_KERNEL_STRIDE_WIDTH_SIZE				4


// Register NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0
#define NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0					32'ha03c
#define NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0_PAD_WIDTH_RANGE			3:0
#define NVDLA_PDP_RDMA_D_POOLING_PADDING_CFG_0_PAD_WIDTH_SIZE				4


// Register NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0					32'ha040
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_RANGE			9:0
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_FIRST_SIZE				10
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_RANGE			19:10
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_LAST_SIZE				10
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_RANGE			29:20
#define NVDLA_PDP_RDMA_D_PARTIAL_WIDTH_IN_0_PARTIAL_WIDTH_IN_MID_SIZE				10


// Register NVDLA_PDP_RDMA_D_PERF_ENABLE_0
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0					32'ha044
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_RANGE			0:0
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_SIZE				1
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_DISABLE			1'h0
#define NVDLA_PDP_RDMA_D_PERF_ENABLE_0_DMA_EN_ENABLE			1'h1


// Register NVDLA_PDP_RDMA_D_PERF_READ_STALL_0
#define NVDLA_PDP_RDMA_D_PERF_READ_STALL_0					32'ha048
#define NVDLA_PDP_RDMA_D_PERF_READ_STALL_0_PERF_READ_STALL_RANGE			31:0
#define NVDLA_PDP_RDMA_D_PERF_READ_STALL_0_PERF_READ_STALL_SIZE				32


// Register NVDLA_PDP_RDMA_D_CYA_0
#define NVDLA_PDP_RDMA_D_CYA_0					32'ha04c
#define NVDLA_PDP_RDMA_D_CYA_0_CYA_RANGE			31:0
#define NVDLA_PDP_RDMA_D_CYA_0_CYA_SIZE				32



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_PDP_RDMA	32'ha000
