`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UWxjbgLc9r/dxO0ey9EVCXWrDRRm0t7uTMOO7aV79OxUPFzmNmFwr5z2vMYcRle1ZJ4gnKJn0Mju
5vVXGJsRXg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b+FkJmx9p9p9Tgt38ZEoaXFBvF5Ev93XCtLuHeoSpFL5mkVzmdXHhbRIU+SC2UZBUQHNmnz3tVKX
KXYpxtwCLl+ozqSuYPoOVpgT7pD/y1kuVt+HKlwAl6Zqgeh+PIGZnADqXd/RaJUxdLE7k5Iotn8f
HBjMEFZ/E0HX+h0Gat4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QUmPuTD2DXWP0Gtfc0X1HucCz6vzmMcTj0BVoEYWWr+iuKkErB2kkR/6wmv4pncABA3w9tbyfs6w
pwnc6yc+kCQs675hCrtprV3Mi77W8hmT8GlfJsibS4C2m8t1s+sKrKcUUbz0M0QfKC3jQgm3RDpo
0ZOlOfJGYL5Oc1mDE/FjrF6be05KtnV/6kpct5WEsw21Ap5T9/RjLNGJzXd+TSv6KTxRPfeOuFu9
AmX/3l/J9jHtpntC+WH7m2Wc6deMIRcIwpcZ92MtyWJfa8Kf7OdA/lmXFwyL0YrUkkZESdHs3Pyn
IPbqjB5JOsR2G7kdHGcKT9AEnfLDPsje0ltRrQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Of+1ixcJtVgLApngBwY5l90wIu4wcE4oHreuLX2dFnYgjXvnV2F2VUMUtvEiwd8rf75m6hQbW0eI
XEiPDJRiJN84rpXLnPGXPOnS3OwfuqRxpFI7T83vyr+754FnwRNhqWghKXD+l0NVl4RDVvQBGx99
D//DMq5+pwS+onntrg3cSS77gamprKbQ0aSxfgxSD42FsQ6QgofKbOxMe4f5ZEpkWraWaE76SBHm
D3u6CDe/OT2Xb22KPrUR8es2cwHVjwQvr6+22cTjyOv+5s5cpwxuGO8r9ikYLOgpwWANipu/auLW
y5LLccLBn4ABxFGuTLc2a/HlJD0i8H6lRx43LA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j58hnMd5Xoy4OYAQg4uUBut8luz3JbRUW3LUIpyc7hV23DnmJMeQW2nryR1ykup8De8v25ecLSyD
23Px88+x+LXTjO6ECXH6GL06MZVDLIB0Bj6943fOhrUhoxLU+rMfMPOd2WL5r33YZt1RieyaPAR5
zdm8bNTRRQ6BFuUsYUVD4Ns3KHTjwLOuXLgXFuU1/EsFMuGpHqfFs6EWzO7nxub29hFHzVELJyU7
JunJhAYsRRJUWIE6HLxaAr38xWmu99OpTb/6KoUiLOY4IQ8VD1L51JMkWMyw1hA9zKKXJ8+wlCJK
BaxtOSerEpxjad6pXB8mQL1wGTK110wW6IOh7w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UxmonX64sEWLBN+yMb418WON/CcRJ7ov0IdQBJ/Pl0Vz6dHskBVEjk1ArCYjoqMbT07bpIlTnsck
/8ntS0Jh3WO6EcNvyxslYf+nXWiWHqNFPTjW5XUxIvxexyOtL6pX1mI7lZVoFsCJs+aC/qc6+CFf
zBxTdN/qH5ETJZ4HnYo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nqWFywteazZhJ1QVp6wwNkFWDAfdm168Egko+3pBXO4o2qRUrrD+7zC1l/Xi7wqJ+X4ZfZk2e4W0
cBzqLf/22uZpTH567Iul7COIsK046KQpVSi+HQmHJ4SYQTFKt8vPapnZFxEqNb0cFKA5BcIuN1W7
YyFA40ArmfYlFjK4uh7pwTvcefLzNdbPaJPhekIZZcxaAJTmHqQFSACK1gmcDcq3HC25mbSQVczD
3YiqFYP1rq6IGerqy3ATxRDvJ2mqQd1w6T8s7aIKj00sV361yI1Dapm1LXTi47jHrBCdBxa8C/WV
eLVO9O+jYuesLWtMjm3azrCM+bFlVCHgQ+cfkw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tNeblXhqo3QnBTLYPujRWZtuHYxesu1bNEQzc9/wNpUKkZg2F1IZqz3dCHvRm2UH1QiTyjOxyFp9
mlDzG9I3JB1+z9KUcnuFtTXikIFjfZFNu19pReZQIuoWAo+Qh/Z+hwCpN+5nkBdJpG2W6CB6Y/bK
f+KGrRv4B0NvEGcrKrbnwwtFVs/9DZSxhYRAhgBZn9vBRsi1ZtlERTVj4LuSjEIPMAK2f1YvkGbL
atAB5GPiCLdc90vIso0yeRzTOs2FvwEH3KDj1/sSytol11uFrgCZQV7HLslO6Sc/EJo9ErT0B21A
6JkecL5liGkXnKQfpdw8ek8iQ03N03zq874igA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55552)
`protect data_block
/gjohAtE18HnhfXFjdgCJDDLircv1wVnRRq9wMXBeKayopo3DxnPCGoOJNR/5CID1tPYY7hv8qnx
0psrLL7LzwgA2C8/AuR7mSzOdfHnkriTpEnVQZliuSWRiNM8NuiRGLMGPiMvO5+GueWtQZapswNx
M+jQw43dFF0f1++nff5+FiZETZUf5tX4OjiO08BP19LNtg8IlTTkxXpbxUiIUZSQZGtZsyhjDxrf
IZBZrja6wM4KbFigBDsSeEV0ErYq6kT8FgsfoJQ/FHQdiPLHQpzH326HagYpTEAPFJ8UIFyFF9Sx
wbOnRby9IUoXDjIMh8Yc9r+TV9XtkpQX0Suv+IeHp6m+e+ECZZCDmjAre2iKHaQ6GBhjz3ZPE5SJ
zWjRqXWqzqiHFTHZ70ffoKOMdMc2tW5Kuk4UqRv/cuQ7zoSbjIhQ1iPklC4qFlbRG9W4zhd8Ygc8
Xk6q/btMregXzDcmWuiEP1eoZEkBEcH/XzQ8KYhnbLyIM1Z3V1TFG0PJuOcgTeYrRh4NujdjZxXU
aySxUeeXXX4n2YKNCaDvLiTCBnis+Rf/xVOB6M1CFLlRBY13CXQpGR1g4hqGy36eVo+GOK/z1UvD
c9iiSQXUcrvrXd6CQRXLi2XV7WGGoQk5xDFjMT+Wyo8RuQJCLy0kDbCWfQrvmSPY+Bl6Oxp7Px+A
3TWXQZui4U0lYzMYuJEeJe8+70EhLyPCpNELkisgLZ1sW5pHSiV9e+JADIF7ffPVvL1QUlwXS83u
TVeFn+MPcRbJudmUxGqSEiopRi+/bHfpfuWNEhAYsF5iC98SUEJQQij+90Mk7edtrfLyhbmTkw+N
YrI4qib/V50bf6i56PJ0DCF9DkvW3/sSUf55YZgraI3k/uH903bCKBQo3UkanVXQoj0DqN/7meUi
oQtHaMWmzqx5z5nJ4Iv8Tgw3kZbrEgI8ybiJoFdK7PFpgnZ7X5elEEjYbxKguTx48sliQVsE4CyB
zDWIX30zeL9Z3AdutiawPPQyfVgRtg4VKi7XbywdhE1dB6HlUr7z4ZKw9Qrj4tdVvODSKNNu9jSa
xG70P2FV5rdf2oRXupWXDaFmLneC2apgtfS1WhyuFtjmBAxyvQ5kVWiZXyuBHjoFucEmiBoQepIN
edaCgbHFlP/NkvK1qw068iqYrHDJdzeJgVTqtK/QiWfOMQaYil4F2zOVhdPoG70XlJCqTa8jpqJW
j+NgEMKdhiGq06Q0KbG4LHAKYCbiVgpnTX0GruOv6MqBt2UDwDUpC2ECJcaS6c9rQ+5r1SD3ynBY
LTOwIvupNq/YvHLw4OKzFsklm6OSJoqgAyjFgG+zAfQ6WeMXmIAAwQ9fmC3ohat12Vtu3j9lrWKj
jnWmH9Li/wxGgxMcrC9py+8xqRkZHT1/ltUy4FcD06Zu1dKOdCSI4bNfDXfIncg2RJLMOVGX+fWP
uDW2YgoYjUWytNJbVZDjxXOqPrkO1iimv8Hv1LMDMN2u+QAilqERzLrRzrUfhDHVP+MAV6N9lG3U
QqS9GdtJuyf//GsPsdlY4LwNubVaQgvYQuSkHODU3JI91NWUKkgFp8xrXfXnqDCRtAovwdfW3Xhg
SS9fPVASetOqJYFpBr4BEfpFAeRZtFkxlRLFll2g1XyLGjNN++vYEJw14Byt+Cdj/dzUnKvmoS2n
uaeY+Td0QsyT4oE7widc+2YatCNKF164TC7nR9IWKjVG2IAKHP5RotEgHeyG2mYyJ0HwNhm3F6Ur
AM4F5ITfhcmAbEwBbf2TdkfBJSxtqX50WLi1q0tkFT2eJ0fcWpATzASFC0hK6kzfZPa7h7FyanlU
ndd9n6SaiZYmFkEOUiI6cOANOClIWhyUgd8ZDsQYT5VK74qfbb+u7/h1ceXo1bgR+sMC8SA6bW4p
IOVH7yxjqci3yrWwGQBkcPU6PKrUXSTGY+qLpqEYrPN6Q2nLk8SUaDetCsH+tnRU1i9fO75Kmphr
MwJaKr1Z4G8fIfbnY5HAmPSdfF4Bda4WeufeUFcQMyG4wJB8LQVpMy1sG7t7SgNYNn71hYhebdDG
cJG5CY4WjTHXcn+1KPEtnpeilwqFbgt7buxftisL0XGYl9LrGbhFVTPNPkDvWfBtKwgdw3TEQaXe
Zi7elGNJfR9boZUVEgSh9xfvL2PMaij/WDwD3T7jj3m6TJhCxOv9xxj7niRYJcg/D37lW4vpliGH
Y1jtleH9XCKGdD5/zN3ikPNrksqwzChBkcIVZuZGKVCWZp/XRzYJ2w2SZWjOuyK0G2z/7dk63qgw
piyf7/JnoYGo4wK2Hm90BtJEmQTmazYhv/yI8UBbbmXd4FEG9e/NdmEiZ0V25cXgSF18adnL0AX6
C+mSlKU2krpZbRJUD0ULxTyGEl8pDKH40u1ZSZ8IKz49+oFGnsOmrHZrfKHMTQsgIbOhw24wM9kl
38THUqtvuvSzIrhaNw6wlh12ylm3fY0YNTIdtlBGT5H0lbTsgpbAAKvZ9uGtgeGHbSryS1lUZ/hD
69BruQ4YwaUWdko4SVsLMktXG1C2AdhajjIO3ZYTadCgnDLTuWSkL5Q8C6PX18XKxYpH1TdXvlHJ
w6pXjUSorhsBp3biN2gAk2LOfBW8Rx5d3LZSa2b+Pt4F/ZbShUe1ozjPBGxfJodvQcxJBZJ34EXt
PTndv4iTappTzLXNUw7XdOx18bbpYDc/0NaUR+HhyiYBZ0Hg17lKUkacXtOzz8VGP7q4denMH+l3
npKYz2gOuspBtJZfcwmTLwLD93L0S30CGbXSxl7SrDSEPg/cbkMCb9BBOutoHXcnzvi1jZNJWis3
t9wRjf8pY5UmEvoaovnX14ypAcf4MTaVCElGs2H5//p6hVCdSl/lAusNTfG4cBtGT4bQkmbmEgr1
0bdJJ2OCO4okLNS+jKjV99vg4ezuuCnw3BFlunf3xRXDP1ozfygpBwqfHz6RsdmS4Gg1C/W8boMx
gmoMHRD8YtITFMGcrkV1vD1mxVDMS6mC0jajplXneLRIWClj+5qyWQPUI/rEAPGXAVUzxqqEUlxW
qMSLvQmnnpkZ+kdCymODvdqUpPX9dHlxLizwEnV2jmNvt7Q/1lb9RS5HJxWWKOFItRsQ+5X5tUME
2xz12pmYCkuFnv7bNDr1BBJHXpVkZTQb5q220rCEwIMNdP3m18HGjKtdRwDWsX6o9B/GhszJz0yh
/Wr9dHdSjJPE9+hDThwFlbTKIZeW/105r2eKYrtMXAs84SLH3xi6OKInNktmPYcRQkxzRBt/0BzN
Vzoc68leaCJZC1XYfu6qsX2n5bXfi9qnuYw6nfV5cEF4MUGMHQ+006VHKABBhYaqInPm/+iIePq0
GNrNM6b1fsXQugMs34Dm6RzmumeB0JA7XlkOOz8rmYUh3ib2QUK0FDm+XLOm3muy25SGHbXzAPsZ
aeZaQvsf6mLXWq6r+Cv8TQIICoU292B6frh6NLJrNi7Pe9k9MKVP0R4MhQblexLhfWH9IqMSBOtv
svDmrflU0PyGBuOd/sEahgfwKbsB4Oyy+kgIWhMwJWzmHEAZFwzoz7NzlvUH+7CCMCbnu75KsA9o
y2OII9e7UQ4OwVTCrCBrnb/LBHxjxfvYGxEboqzrioLXGJN9oWNv9Cor+KygsMM5lWwJok0zFh7v
XD+1ETyx7c6rP5jBIeXEHV1F54e4a+S4HCOwFV/j9S3bkoo5AVbBC7Im7wpWCBBBSAKFzZ2bJPmj
RVp/wHVd8iNJn9sdUWjVbPzOgI9EeUZrDN0G/YC4gCFd52xy6IcWPVFwWGvgEIMNT82UKwQoo8qh
ELZaH2zsnmDvMUwMXyiT8QmaaOW94LLicqxTejzUJ+6H/2gGgU+pA2QaSfoFlzuYW1BZwVCR7CCX
9RvmY9DE8SlsQJouqJfQQbzoKCF504M54zs50/ehOdqlAcl5gNis9x+/OYkGuQBBbdYofkbiMMwk
fp1zP4RoEIGIRDxHviQj0slQULgImLLFhLQtHrVZiOrzE09VSevGDN6b3+wJm1THpoJWBPvVR2cN
VaIEbjBQy7cpTMn+J95psCCUxFryn/Nr/n24LfFSmuAUGckofq4Rplrzg9LYwzxbd5UeBYVqL3Q5
YHDQe/g7vVFOiHUGWD+SthlJJx5FuhRySCcb+w8BhrNbFp38xI2XB/i4Oj5mMUAgcy71DQTUIZYI
p+GHcux39A5s94roxGvnz98QFuCF1yrLC7QR/aUMj3H/bPKgbC45MSii81z5NZ986PtLqX48+D6g
dxU96baElJRoEdvpnPqiis2c/na0dv1mPsYdrVtLsr4d1z+BsNPKph4blD0887yLbuGjYNtwnKA0
sWXYXqhsZeKHcgbpEkolloYVNht21g8wsouoe7kjeBtD4KNB7KiMPFWOxFyxOBlL+E0BCeEldE8c
QRBPeuAwGPviqhHV8MmYJagM0bvWbhMM77BgZ3Zfz4TbBN0Y1GhW185GGEiEhI4W2pQrVe6uXp3j
y4JQ1gnWmTW4rjCj5zrlMdTfZN8Vk4YZeIVTpzYiNUYTkqbNEEPPKYx8Um3vTaIaFvh+XFZqb5/L
1kUiyIPl7krCayXtbfFuEJbj7mZVmxKXzmP2fhLBJJphe6LBK7Q3WCJwTX/Ja3H5KwGn9MWFcw1O
p8SZ2bljcFpl5Yeq86JYarKAW1Ihl5zuv8QaIEaPzEnj2SQMjrkfD5sysbUhf06CXwFDakulasZw
qUKwaHZCpWa4cM2k/VanLtqD6qqfbxG5ZNqhO2ii4LAl1tKkmDc8bFRRnJ6zMxT4/EXJ+TK9gkjM
b3FrMXzr8e36VWNFtPJJoc3BuHdN9gmR4l6XQ/eytGDV3jry4JSQ3DuXb7LR4e/jHvLtw1kPz3hB
4pN/WZxV8UQw7xao+aLAUtVc9UWCxOfJxngX1GG2NbcITYKRIhlVwW2dwCaDj43H6CskpMMmntho
OIhOpKuMwZxGswQ1X0TP+FKKOJ5Z0ObztEzsw0ZqHlPQbZfsTtYGaSTHRxjvmIBhMMO9iToKjv5P
bL4g3pmvHaH5ZTc+K+9R5Y7cUHvzFf+awAaU7bKpMVmqEFYF9/RySynyxwOHLhpd9hVxdadnEDAX
FdsgBXxAWrp7f18swjsm//+jMPiNoy5CF5HWlZxEoMiaw9M9Y/uyW6nkEi5oWsJSInWmq6RBGmNt
J3XGOgHoPrPSa7yyf8xmTxv13GIxfXE9LcbIwPfSwrV6MEfUnupeZzIQMlfYEXjII8rhdjfHepa5
DJmbXLYWDooHaPGeUuzRCH51zlAJrApR6skKanDLx8J4KKHrNxChcS5Clxc0lXt3QlNQGq/Obybk
a/yMUASkRLZ97UiyL7n+Bj4/Puxjk7x7RrDuMckOnrg2t7HlgASEQrqLuZWhRAsTAVw8M8x9nLGB
+SGgFwN3Q8QNMMDYMYMNS5Dz/MMx7SucM4RonPmU1O/9Q+SrMevS2EZ7WAqVKkvpU1nYCo1sCuHC
XMs0Z1b8LSCuT/IRIcg6xB/fpZTVDxFeTkSHsJKL8kv/xmnw4ysPsoDaY4pdxvHF6G6IjbcJ/CQQ
K+Odk2hKIwNxdNLSiEsBDSXSIURhb4ZCF8cA17HOgAaZ6zilDmiTGzpwdZ8KSrnUw2EbkcH9my4W
tbh+2iAaAgZoybNvcs1h74Heg974lXnylc0nfgpApbMrrBO35Mv2Bb1VbkGYLpVzF0CAyPiGKsep
z9OXOqRmXQtOAHnHw/kHBECVZILN4G9rcnbupq9aT5/+DB+8/VM/wvg7aKEJktlDfDhBzQDIdR/1
iMA5ndbhXv63PH/q5JGJzIUP3Q+QhHcQi+8lK9r06MuAFoTkbE9xSQTNY5q9lvEb9w5xJlCGziDl
5QkdJ3pmkzLLJ6QOANv0lGvzh4khUz1qZfv0PnuF+UPVEMpamk8nj/kaxfDz9HiHHwFAKgjm48oF
zZC5k4oqOrHPfvRnJ17dK7ym32WaWVhWIUWH6lTvR5RWjc+GGOs82HjQn8XegGeWyzSjU/wmDVTq
zRxCWLSilUV013JUCtJTqXqOF3FgWmJd1hfx1cCSopl/Pn++mANz4FTdeQR6ALSgvb0rHa5ZefuI
BLWOgX5RdW0rcWRalPvRkTJ5gu1pVlRRUcr+BFNuhLV4lWUsbSsgIOT3Nm/UhRmroQWKYyQYbi6c
6BU8epjz2DPSQeZgNQJ+3QL6qVZnEfO5qGSyPmmKx8dikzVm02dw3JG90e5ZuLWpXWZind9agB/1
qiOk+SqgkOFoH+lZwLBqoL/OcRZLwxF9FPYa26D4MLD5z3HM/4wjMjtkw2xFmAitQr+OKqfBIBi0
sA+XK5gS9bAsYt+Vurxd78un2f7qkYE53kN79V4t8L2vgdjGvAQFa9U0JaLcmzmz7EGwfVrtSQLX
JK5rPeDUZe7EAVQzINncKayBwY3BGbfPEa95l7wEwDdtk9NppOdXlNg3imLBxNPeOwQyrKYqR7ua
6UNYr3DavxfFbwftp5gsX5BDqLlt6qi/dirzFXaK5CFkc7bqTnr3s7KqR2o71RFg0SyyajXlXZ65
dJe4miJEbMurlfWCHCzIlGxYYiRFV5QEmaBjHVC4jqw9CHmheQmpoKKNJ1iWu5R9sXbCuWqWXFU4
E46hxhX3dykel+Pq9cUV0Ozu1mZiaOlwLBUewTdKYOcvpqE7G3QXTXauhkEhUy/Tti4oflvmDjAR
vZLKNOOTqujQjONiVY7EUsKKXH5M3kwPiiKpGb/rDX8CqyP7EhjAALcPCgEvftbWbyJhHhIdVt7v
opUE14TpjmIIv/wyBqiFJpXJW3aA7aDzcNuWfOu0ozpMM1Lg1myWNADQ/AZcmwIcgeYaN2yDzjLs
+7QmZGZh039ni55jz7d9tqzDTCIjLy8QmSQM2ockiV63E3OfSM3n/ZQbyJnpOxWI1PwMSfg4P4u0
Kr38v6cLBnyzZ4GTU5hcYbcPcJ2ZILMNJi3JF9zAftzSVoJscqDcNFBHY8mL4KAq6uyCYCGaKaIm
W2vCdIhxNtIkAuiOwjVshp2Gem5ypeOoueJPqhziKt9U6v+VWisVFyWnH3BWshZxl8gdQn7D8LtY
Ba1vfjp+FfuQgKLWXL6MTCun3EDG0B4BZ5860NvzJySDr5BkbjWPZmK9gonTZg9/Bnx/qPYyI0md
hXdpthhRyYuX242rfxvmFMqJCONuHVNYC2ah0mqpKh1W4z4DrLuO8V9/N068Ikcdg+rOTzK2Ly+T
DZlqEEYn9YqDrZdLNK7KGF4OU1MYVuvtmRDVvg6Fop3TM8+pmi2UdEt6zrHOxRWCFXTx1tEvfof5
ufqz6zR5ls+Rfbg+xJcDcOKu7TlmPE5Q3WZsqvpwOfEfgE3HrlrdaTOtNTdKceAG/GLaeovefcQk
4UvGXW9J0M1LwlK2PvXtHAjKhm8QdBl/SRxfRDfReX6yilD5zGptE5EJLjgOZ6Pi3W6bawNUfzVz
uaNri2Pbae/AocMXdBbNLkHTYN2w5DNPglWUXuQPDEK6vGBI+9baSdoYr5s78iPDidaZ/lok9zWC
aiOVLUnxwz9qOu0DND2sEJdPrgJHysHvSyPstlIWwpN2JJzW1mAFP4HEfdWv1Ih35mNX4UoZBg5f
zoboWRRPMRVutFivBZgPh3ylWJfxsVO6ORVyVCwyJ4NQ+ottZrNSNEJtwkRXZlNJwwW5sK0eCbRd
WedfHIIpaMXrq01pT5nzXTGyUH/UsFFscwxjksKYNeWedbHYi9Wjy3LIKu6jvmNb+NImVzgcO1Bn
NNalueTRZTnumybvaC+98/CeoCH4DedMmlcEL5/79S7xbP8KYKqH0rCF9ikb3jnnj5UYrRDeWMfj
OTxJS4yBMq9qRJ3Xsmc7HSONdBUS1MhXiuuVJ2BA1O/q4G0GqpDhDTA2uvfKwg1WopAyPYy/8Era
yVOHfKQVWmXEU3ItopTm7cjJNwUiRHfqIefl2nLJxV8S1ZjMNXGRQ7N2ifTZIcwIuP39zHIkSAKw
SdHRJS4CD1no5yWoC42d4SWbf2wEY2P8PyB3n+Bhusfz4lfNe4k60Dysdk2U1j6GygZk4pLfKEjA
4TLzJ8pwHfi1J1lnt2dDUuhA8OssCAWxjFFmvMbo4nJu1SiWYKMpTngnYRUFzwJC8HDcc+zFiJh4
eCttHAyxdTssUXi9pTibMrEL1nCadrA9kW2dRucmCqWxi7CevRP+lbb3kO4IIIWFBYi4Fe61R7ok
83HEYgHECrgUECzl53HUYjbCMILrkIMMp6EMlHcCuoeHGYZ1EDcsLdmL+4+/Rdoh9NpL/WXut8J4
QxS8JhsE5+cJJZU6XV1PHgxCGiXN/DuBErW45HGzlEHp96F6M2BJ3h4lNmpfm//DpslfRh8FJoaJ
nd9wJZXq6jPWWMcAGPxTyUEaVQwwwmXYeypvf9N3Nbjt06Wl9p4Izsom2bPYdJVuHiXNpT2fAehT
G0xJhsM25ysCC8bCLtimZgezxxLIXSkAFKbcV7o2VxxapEp9djF60JzypvnChefzF8+9FFPWJZgL
KXFCKo9q9RI5AexBJRugquwBx3AtvYrTeLVMYaqocqMNzz9Uc0Ira0wgiPHH1Wv4EHhG9LuDUcqT
H6UexG8aWinoLKzmTitadz+XaB1eZoD22IIYfNQVBwKq6gQCzG0oYy7ppOKPvAhF+4SUUb+QTUal
fkMeGXIZMxGxQtMWzS82k0IO2M7fPTwI+bQcEVDacnc5x9gwBPDm2o4FLZbZ5ugatasOBX8NFTaf
fh6gR3HY13Lon+gkIeQprrxNmpxVjgbV13DQDhTEmoyKMIaoIMKTCEDZXVMRuf1u4ZRq0HvenFAQ
A3jngaIHo9JVvocLjUwFcsIwMqL0DzZcxiqry3BGmjyIn9H40bewZbjpdFRHFmUFcI10smGh4cSo
a3gkBKeL/G9XsXfHUTaTuGjjyuBu4ps5/m0KvBoy/U52eY4Fv415jxywrGlyiTPwIN10Qh0Gm0JJ
BJp+8D1KmEXDjEXEUzJ+EGBJKi11GypOFXqg3x5yKv6Ss/7yVl982v/8pdujWBTy4oi/95DZeuw1
raWbYszwfsjIH0W6lMokpBSa6Im1rbNz20hRJ1aVHs6EMI1Plct0F0lDGP2fwJrkFdkAzSPSSX//
fJKbvKz2w6U2uelZHT9zblHqL7FD9vk2CHTcHZMrkY9pq5//6BsS6RMd8uFjFI9PQdj4ONBqaBb/
NRpP++q4FXQv43vzQfHZGM+XGjwNwP3S2yr1wfD8hbPcvKwjgWbTqWpWYmpiempwVAB9CqhLB9Pt
uivmOTW5zeIpm+3DXF6URmi3wXL0QWVIEuCnKTgWN54cI5Ayfz2OCk9llA9LJ4ixsS5pDut66g0v
MVwknGDsSny4BQjTKaF+hc7ei2YiGV/YK2VadTQ+2U+Icw4kV2EdufT5g0NCZayz8lXS75SbAzLE
JnPnjfWfiSqXRE1ArP6iJEhI9BvP88pdhwSey7Zq7ThJWl9rbOKoWRi0TaBtgQbdbcsqEafp9r1d
oynLRN7USkgLcAuSPV1dGhq/IY5Mrd6CF3ZBCFBCHzlFDauKvGLqJBlGKKmJv/t8mgnBhZswiE16
Nt1L9YysYKujxY+niaOt0JE3r93uU8bkkzZQFAF4U/qdvlaVwREIVS/E2Rh8iZpK6L1SCi1J17sF
mrOze7MoMHTBQSGIweks+2wLGPYOQt1u9n6yHH59bUSWkBUwEe4Z0Vd58evE7uolJYuEvd5zQ5YB
ngiiHor5GiiG5CMBMUviD21m28X6Jxs5pfk/aUzUOFv2386NF9QjevXVzOnZn3hkMysh5CWHsE1K
sIp23rCt6ozCdxSocLolg78Qk/Xo4pnAxxzPyCFASCl7lUgwjqL3veAGOmDi/4m1gXMPADVdi3zq
tk9Gt9/K8z+iq4SdSXOS9otnsQ/zxZGMjBgVFFy0kHN3+J5VMgvP/d7/7ACdeLJIOHF3u+47i6cH
kBlZvhOpQEaqBxARH8JTfgc+hRXa6e+b7XmKRKUO2rca9isrtF1lhBqQscHofYtc4E9cUESV3SI1
eZ9q50x604swnv+KmJ9twBh/3KUxIw3ShsrvydOnx/zm9BP9ug4u5mTEnBypeIdEKZgpK0g7BfYM
Yk8F0Hjpy7ylwi/sjN5G0N/1P/cL/V/dWsZMvYivHYXBl+/6ELxfPz1PBo4nsJs8yD1vt5twBOoO
yoDs6ihToonwBWaJa0BQd2FinFv+zEpWCEDa2aOYBZ2qS5LG445qopEkzuTM5hPy3ufpivUvvxf1
pN9l2JqLtMigds07kxCPQcvOlYRCwv/fxQUa8UjW8lTpxR4HDZkOq89Pquy/h/27B41gvE+PAxw7
+48Eg12X0KRfzxs7kCHenkfAwQSMpMuhQIK0CAA3KDWnH2jto24PniF2SN7/mnEUSmWI4RQE/zbH
0C6RIjVQg+mQsFjxoUo+je/LyjEyq7PhFo69f4luUCqt1qqnuAgk1H/mIdDb2YSDnzeGG10Wdm58
lrQqvuw226cxhVxuXzQn8lUSlBuRCxI+VfAlRQO9+R579LAA0tTonERdfy39i2MODlFiQ06VMw1E
oidlMWrmYrO7anroyxP0G4MOcUelk6JM4BgburlO3O3qIDOs8utmpOLPavLB0FKJqUQJ2covIo27
aVUr6LyrJeuOMi+riI1+nvl628OZLmJ2nGLac0xcgT3fVRjiQeOkohTxGREch97XP54a5so30+l1
AaT19Tk+Snh6hS/atDmSIQcAQsyvz61KJgKWmERSJ3sfa6zPZYg2NTYb6lCaIwjxPI6RSp2QczkR
Q+uVJ5pMueqdDyG+4EJC2tbydIf20Dfep5/3OPk2ujn6swn3TNjMIRdgbLIWP+/nsdTi4m8vNTfR
Mat3htC+UGKD/UuNSuaHbAP85KLp6jjipRcGRwuSKukVHkNRSXrfMgmcJmcQQw6l5pFojyFkymIY
rp1V5PhTflpnxsUvz8TvZrJ7vTOWLZUNfdhPiuwmqv/TjTy2AXJIvh1ECmD0uGSlRvZ/GCKg5oBk
doKOUeOE+iAgMN6U3SL6HhmVz2h//B4p7wa50xoonWEFiX8XMbuNoYpgMG0Ie7/KTToPb1TWJIT+
D1qRH6insTABItbgR5UlZZCe7IYOAJMvsno+5YPwZn8OihhCh/7jKjFYsU7Sx24yWCdZ+TnRUT98
rkacD863JiNoGgnlZajynD+z7FhkE8ziPO2795fCcf89a8Y4jmacaX8rJwn7MmhQsUoeVwnasc6O
5/OKM+sNj+dvSHtspMLoMOQRWxp9jQDZYOUOmvWhoa7Gw1PEe7uf8mb+2xLoO9ILATg1HN0e0W9w
g7TUq/z0YYjMiv9Sa2LJ3uDMoNOqzmZn8L1Ft991Wzq/KCQ6QrJZUQ2Cs8/rrhGfACSnyN5PSWPS
vSn28aQZnEx5B2WGj6A25e45g16ZQrSXHElRUhM1k2EG34w2bmIXA7c+2vtqUoTa2OK5jjv+A4Kp
uupDyTezQBA7agjDlkV6dbQu1eq4hrZQFlGYzjFX0yoGFjEAdV5PoiBExmz7WqEsykHmiwt2xS6F
sUEwzbP+6df0bKgF2P3v6hgSceTHdG8ueERUxuEh15UDKb/jy87J54KOJqrTnq9M3/i15FKpbL3n
pn0/9l/8N/LbsNct6n2QsoNNUEuJdHVt1wO2Hut3x8v+7pXWA3LOQBJ/b31o47J9suTvGhOjgs1O
5q28F5+paykCGavJw4nHwZef5dD4yIM+saRrtodaemo68XLeDlNoaSRXJTpADOxHvf7zHXJunsYv
wOvT+2afyRzkzZqa34G+tarjbUZW3gm0PRjUbMADD3foUBitTL7ZLIwMm0SarDwZkOG/Ph+8EFAG
EP0Q7lnslRmpJDra2ygRgii7XDhz4BUtsXE+cDmbm+xucHneGxakcuyNIuBXjlyuv1tT5LBuuZyA
BkW+JlnBtFw0bz3XTZaQMw9ZenCxvYHS9smMBqIwklhc+y6mYAqk75oiLrHko643jwQhQnd9aZe8
akQjAhLMGs64Ccxfjndmm9X3oM0aeLWcdgTXmvfjkPMIY4Fq1uS6d99Y2dZsY+OfDgCmiifzhzCI
TgdQ3ezRj2sPSL0xRCS/KMSgEyrxeBAo3Ltiup02uEx9oNv83/j38YywHVg954nZLbbT+T1Mo45y
ATowjOUXv64Okuyy/6mA7ErYaw0IxXBtAfPL7GA1h6kPK+VEkOYIY4zFLTqTve8cXqnOPocWBPSr
zfwIJ/1rqKgjLZ/ywcpm0cFh+CzYpLYzrwr5R0E5YGmTrO7Q+9oaMw00QUmstWsMoFMs8eh4lZ1Q
00hZAIuolNefPbHPlHhRc9Raaprdd0xso5BERCkeVRjE0RRcPYNYp3Uno5sDQppFssZwM6HwxHHC
8SX8hyDNp3PprnFQnOE5CionSK/U4F+09trVLXyIvgiw6+ra7lt94yn+Y1IuIexwLLjLfMocQHHL
hEx0akV50QpCEx/wiwDeapFoeGEeClkO6KU89Lyq5Ol5AYAxe8ahr5EdKECNyAe3LuLhufJBcoOX
mKL+Iiq0LuXQFkEYhD86fgI7q0ybQeljkD4rssBHN6W3ALhNgEuiK84fSXLOrfnpxdGgK7ygnIdr
pg5UzUcMNlXK9uxGq7taTlBbEgRfbd5nEuyOKYoRRJARc6C8emu9rFkSRf162RZ+smNLOp74CnkH
ncYE9tvIYDsdoas5SCRyACi7iZMfuRLgrsoI/rrpFIOML0bR0hDjzYayXRuMtveWudJPJXawk12m
TPAfibueNDbOw1l39pyZMOg3uGDdb95/d69MVBtFRXDMQj4JmNZFFEiVwfp6i72oWNVsAaf/gJk+
0jggzYsDNzPSyWdzjuh74KkoCXrcgRsXR/FageKXBbviKE3Z7cHIOZUaKIYCClNv02tCeKUniBnD
4BR90IegpRhlDvDNxtRKQcUJgQSC8ywS7vr364+GWtjvpn0yYAQSfcpQwxsv+vzuKy5x8Jdi63Rj
afZsucI62JZNCARcrw/JAc5hTsMxqPVr0v4TG0ioUPuA4p6dTae4b6P3Qn+6/g+AE0IiC9k4JlBf
76pMEsIqP+fO+X3DMoC+9xp7d334lpQcVOdZQv/Ni1ylxidq35Sp2C8t3rct3FCAxhKzj6ThZMXq
vLFu3g++cIgKB/zIxtm+gHxlQjAit0L7UM4tnBlOyxXKMPB8rHHw+DJoKUwKwuReMO0utmqKLBfs
4y/3RPF/oug1gyu3XH44OOH8wk3SLjMiO+xuF8c3nZzB4BqgAhpuvarAlwM0u+Shcx+2C50NDBel
4TDtZSIEq7bKawjaIWYzOHagdd9pnKEZ7wmN40t/4b6e4TuFzukrNB1tT+b29PWM4ecyBB4r4eS+
fHsoVf0zbqQU3nWc5BzstCw9sjshWNztmkoPmTIlkZeqBiQJLrORUBFtogB+XRumLtHPm0ms6kiF
+3Qc+7xUZkwVmblixSDZhbLW8R+umF9QhOGddBWCTfzF7B125NpzVqNjazGa9hZBjl1oKlgXevcz
wvFdJ4ZTfYXbifAOw1A/YMCJIfUaNKp4ivoYuzfdW3Llvn+7qo8kTm8LIUN8MYVXGoCqtCRHhI3d
t0jh958XUUDipKeOGpDkdFILf1Pf+4TwJ5PWin217nA4dCP3e+4juQ0T9tM8Mhyd+2jFPF2hxKaM
swyXTVBJAQaqbt/TIB2Z3qoQlRDT+O3GodOYKhByLcH82w5QyKgOp9WORsM+tN/ipprvirtre/zd
xOzQ+K9198HfqSAXvF/zxLMqEO/1RUPTe/tqIT/KdConZUrEDdQn14f3y2xJ3c2MMEaTGqiI71O8
Vt1JDgKUg+YErPbJywFAHpE0InrzE8dDPfZjtoffCC2IE1dzP6qFAg1zYAf+LPs2ZAQxQTPuTdfu
E2HUmCmBcmOUdQ6ClM7+whiroaCYauAyHFxtEAjHpx4O8HdzAfRUpYuYGNfuQfBwYWRMuMmo1+qw
77vhKmpd2B39uTkx54SNgVrLNZ1YheygPAP7ABMpKUagZ2+6kJpHPEFc5QKLVLdik9pIuqoy/LzF
sN8yXPevwZNqer9k44bQf9EaTlXV8NVFFGXGc5vSRAvhIUQHWpVkGL7wQhDvrdBWKoPa8S3/vC/M
/51eQAmqSdkwC4qUTylhwko8UEMP/u9IDBSnPAz46LEf28uybEsMAzxR7mZtVUwi5oD9Ed4ANUoo
0l4+9xvO4yxuv0n27Qp5dmCdDpm6b+LiMKcSBT0ESRmBfbiHvLXqx9Mz+P0IpRaOWUzZVhULDibq
CRIPCN840ZgsDZZ7z6bdsgeHmbXRmPRYslHDYAfDDc6GfkiB7kKrMxEpyTs4r1bVmhQTvPyjwwhY
Q6IbwKgBmMWbQNVxSrIErkfvRjuOq2jYGqlDUWXxremkYOK25HJKBRGHJGM96ltEslyG31j/yC+U
mMYL32bAqhZ21P8WoNFHHPSpANVzdIqt13r4pEre5d9VihcyLL/qkkUj0TaA9xhKZlDJWsSNZY3p
dipz6ceicRomhxJu2oeqeXO5unLitaMJdsiV+ngjI6OOYB8IQ96SJ+Ekb74tlJmDty7riJA5UuXi
H38MHKXPicfHqvf4GPns7goq9UHN3Jf/clA+mmfdt58ou+rT3Z2UrRFmi56vCJnOrivH+9ob4S0S
X6jlJBNlRh3PtM2zuBoD58jKsChXUzBCuLOfNKgm0pXlJdDaUSDgwmq7wHHGkRG7bKf78M32ovFl
1pAW+ax6O31JYQRj9eB3fUypuMbscyCUS6XGuzS+IswqKGkibocQqafrlEs4s6dNxSHjvTtri6/L
xl7DG6RwDUASPBWfSJNJgmAJmNQBifpVtIVShzUl6ZxjK3GVRBR7pFdkrEvKNBVDNiat+fbK/Wk2
83+wkmrXg2SfxzkDM5CtwqDBdDLIkForrg9TazUL/PIU5prliiziY4tphguqxtsOmgjh3FlHa/th
a/DofVG1b56oMBGhJ31npYud1aihUkFdwaWXsXbPQ1rfWDFDvj5vl8JpKGujJovyPQU9NSyiyz4I
YWsRu06b8gTOixkcMjJXi3ShV+tdQw+n9qzcHbertmiPYz8/nENyxP6Mb3QN7LDD0UNJbevD7y84
0zWLxGYfP4cU0nsUIlP8WpeWPNs7H9z5aFyQ7fjeyWO7pDHOhZxSfLbtNvQztt9cbT/UHIUxRDzp
gR20++O/2IQXKO6GcTGGHdnpO1xuaNxg9AYoseE7GlJtNJZBgS03s+pEhxROtrIMItdzY8yfPWMG
2QBlvHKeItq/jgDBSj5FfkPPSEo8HDz2+M84Jg+EcgKleV/RZukYFdqqCS6WgsA8EVMFeAN3foIE
W+aaKQTOz3rZIaf+pb7xb3JlhOlazdeD1/PP7GMjumJ2fkRkioLhB0PAH0FmAaurBkPqkh5xFl6B
5XH/Ukmd8XO7xDfjh4nbeZ3vOo4piMTvPudmps8mcF2n72uB8e1y5bOfNB+od7LSSncKytaJKCBO
67fPDvBUa+GWHAP20q1uWrVdFfSgl88eHEHQ9zwiKpcsTOfsWyz5uRptIxtoyN6oRRsK1PNYg7g/
Sq0Kq7/yQKGDiMxOmamVDaBDVPFObhDj+L0s5wcB3jnSgenaC+clR4fwzve7U89LqqxIltx/n/cA
R15Pt65mIl/CaDv6YgJEHmPzIC8dx30qi1LCj5KuWOKs/0qsR7MlJ0NydwEdDS4K5tSRMxFpRoaF
Vo5o4rtL4HLnqzOWGeCboLwTop7jrSSkYNVTPQWCkAhfkvmX4R0ncp/jVM1hSSxju4Dq0RaMf9cF
FlOtGWmNtbRo/h+Vuj/m8DNIVuvecb2KQDlcDV3BlekHA/MBctTSmq6tIuT+j86klmyONfx4CWjT
xmZKr+RqnKwbz2m4/Hep6I4/lbHnvFniiXc+YHQb6H0ziwczqM59FyhnO8NaWZ0m4AoJIG4oLXLM
8sSV8RChf7L+QtPvhKq7gua5Jkoggi8J+A4DmnkHXIfYBL2tLfZIWCTTxNI5tXN+WRw+7Dcth4m4
AThmy1bUexzg45Lnl+fo52VPeNPMryC9GCF8i/gAHQs0/jkwrIN37TfWylgyoV10KE8+T4apnamp
q0utvW9xPNNGFwcOBrRsOz9hPdbEaEtjCHakZ1nn5NFhLi7en8mG81Tru5h8betm4HknwDGDKZFp
aohL5bMMJmpt1T050blvzesQsDmKSiSRpWtLES8e1ep5evP+8sjIJPs5jieYOST+Tfvge8Vuw8RE
xedKSh4bQI2SUHCZ1yycph+eWmsjKO0zyD+wcGwVvun4hPTvtRq0Mce2IGFqEkc8/0k9vD9rLdah
tPOh4XBcrvePuNpX2bOlGG0hDC9hQWggobxdht+twhRz7iZntF1Xt6X5aUAwLhma9PACJQclV6f8
yM3QUeovJP/OSlEl3k1klzuLFuOIKXiCkCeZg5KJRZK8pR+iyEHry6sOBHP5aVuqFD7Npp96uLWU
VQPZUKFKJK+2ELqSkP513P2IYxk7KtZSCwpjOHfgHWvxrmN1ldT6DFgFn5h60hotr8ND5Y4Nwztr
VvVyvhHPzUa1cJNxuNjP7Q4PRaHYeatx5VY8gwHRBVWdyA8Wmf2z9W1KfrrSG6FTPCkIBV6QjKNc
9vr70Py8DGg8JZVM2UzEfBWfetkf4zI1DkcOG5sAQSU5Zr2PA1jIQ5PdHVKyYSP7LVZdMjP460e5
2dL7cIBTAEVCwvQMkx2+bZy85PjhpmndnOIjxkhB9vFIXR72udtDyXgv9Tho86xAJzzT3/IsEWHO
FRDiDNnFtSWD8xStppleYc9L4XbjgcnqiFsPm+CeNsGtzvOKKcPX1rRvpqOlEPiAzFWNUqQBI+Mw
X7JMpbrVZgPNXbxTI82bxVE02wC1XijkvjomZ5bP4RDxCwHFV5WtqggKGMh0B8cD4KIHrfUzM5Tv
1ajVLdsb17w9efLsB8t4dBptBlXlygPcMCKMMts208CktaS1YWeQ+FGFeODaaMpDsQ/J3PTBoLla
x/vwKv8wUzpF67+KNBlhYkqkUuDUsvB+I1ju9WY0fmeSmdWEg4HV5AJGP+JKVIDvLL48v7YDAPAz
syECmqWjC5l9e+TClAaJ/S8nxCgv8S/vzReIDoHzLXO/xYGGx87R/RKPe0+Nki0y3OCVHd5eoZjg
hbE46z+1xR3U38ROTQxIn5IzhomGReDnxl7p6qRMoXTGkD9mDJVpX6rD5HA2yITjDPDm8Xg4kAjj
eRQkG2NtYOw3GcJYc/2m8uDa9S5xGLumsEnlr8qL4xOOHKFJ7ObVhJS6zFtO2ymMSDB0oZj8wees
P7ZDK1qpaef0nIgU90OxufcucP5AhBccxRkZh6RB/JYf29QzhsYuA0Yt6A8aovR4UNu6QEon3OMe
/zi8UQ6VwGOC0NfPLnbdtdAEVIpyW/19YhIkPi6+TzxJx9K8Um4N2Zzd2xKT6rJCBh+Sa1iYLxEd
1ByI3mSwhXuw+L8JV1fNVDJEJ4Ot4UbevNay5KPJKoUp5NNVqoNRlo1dMD6OQnz9Dp87l3mOPO6+
RLf7MEO7zsePAbXkhDHze6KxL3/wmt/fJJD817PqZRs/aaJrtDJl15oPlRjNW7Hgtp8uxXByJqX/
tz59XFe95uhb9/RQBSkyBiF/4wi1Qr+ULMsz1slwxM89DC3DafFy48Zri94WcQ3l89LH2mxCxZ2G
m7XPKdNTLmsYRdAGYUklrYjT4OOucPIvLjyB6tlB0jpxw4ChvJ7xXgNDEc3Gzfrv3UllG9/riPoC
QrC5nmYuop2RykTE1uKUXsOfjS7DfromL3kWwPFNk5BIIyvfJumFijLAUCOTYzD0uMeKUgIaqh1x
vyh0bzec62Mru3fWCQTAONYxcLfHrmtZ4G+R6LKzd+A2CuIJO3Wl0VrZWjigVYH2+o4AsL1nTxwS
vAJswfGDRPRmAMqq93N+MvDszxL6h/5EvuX8b1qzS/NbWIlcRyy+CSfrZ+IvJ7LOl9w2T2tYgHNu
vMjCaLFo3MWnqH2kVvbgQiFytcBUCS10Eu+Un2OjS3kzW25rkPpHl6/8NEn3HmAPuqbIhc02sh1l
QbWZmnpeHcJjn1MTJZXkIF3dw39x8SEWvL2/kmgLI8SdPV29mqB/N/n4fMYYDcAKXnLoJiIcB6eT
Dra9KXReju5/6ZV0Kf6OWDr5pyHSrZrPrY3OfhoRd41NIQsVup/nxUfNKU9faWDZqF+UTG6RJdKf
tq8+FInVeJnAh+wQDsrRKHzlkw4JNscQsUp1BU+4aJQGMDmdcCBTh2DVc78nNzBz+AicwsoKn2Ve
b8tm1WUxWODu/X4Gvphw5vRj8YWl98hPoMX3n+WLTrjvSDtmjBq8myHlr7Z+c4Akc6RJgaFUwebL
+t5UzqKZZ58UeecCEnJPC14guqa52LNgqY3rVJhdhqSsNvOOhdtc+ALKgV4l9QX32U4ARIKGU/Ms
Gj+wv2LL8lXBV+PVUhdfgpiTrUZib4DoPFHn4C7jAklcQ+j8a+FDyXDXvDOjkuLAiMRQuS5VaAjG
sNjjbJBtb7dVoE1aIb492SSbVHpRXXssPtX1T9MM8Ylf8DLx6PvgUdeyntFI3Wt+SBY491oUaB6R
ohyiHi+7vcLFr1PJssd+y5HhnNxO2opP3Fclh07Cy2p6LH60l56H6RxaLMQpkYUT45iVjhrcJPBR
eomhVYjXf4Zo9NL83aEKrEm81APcf8DnV7mcu0Bc+0mRCtp/rKYb7LHLbizWatIEm3nqD8Xlqp6J
tEg5BM1Kwlj0EEPzjrNjSFWX2koTXwIiWcj/KZUHIVRV6FnQkOIKad86cAdgpen8/yHziqMHDlMg
72etPs+l70pmyK/3D75jhvVpyXw6l7fEXQt+Gm8yTvQ1j6uDQ/0sR9dtUZOvOwoTZ0/QWUtm5N70
KbxpPD9dL/fFYaHkRIFspL1eXY9L+VoSUKG7RtpNZGFch1spYjevsZkwzQGX/gaUOmJ4qO6Vp3rr
oyogmSqOuCGlHQI1e8NZL5D4Tg/cL78Zh/cH4tiosbh0YvvKk7fUuU4wzdu19keRuvqU6MB24DQJ
sCF/yRkb5Bjbu+UquV/bpvHGSEQsD7PYQDxrMImUgctIimVqlb84jpDp87z7OcEqqHyb4QCkJ5mQ
ZClmFdCZ+bwAILhHtQ9sGO+QuTKczn+9VUeryugIla2tWn7ac+40oyezGYQjcvUEwQegX9K/88Cs
mdBP0EMMZhLida+QCUxPYACudiajD/ItvSwp+VloAlD/uk8cp8nZZ8hVn1B7kyTClWV8YQ6W2Rt2
Ln0zfX/8F8iktsEVikyjFrOe2A2ACGB9+Hx21qTJ21+pRR3i4nqqvGO9QMviqZUfAzazhdTbu25R
k0Dvi7QRYLlxVzf4LEd/9AQ6tSkua1i280I0seEW5KsZQtSVNollLt5q70ylWzrQwWy5E9gw0vIx
g/KhIFbu5nIrap1V3g3TVSe2yYvhXrNv6d9EOL3er0I8a5WzbHTVr56dhPOaJSxjxzekIhiOGRUH
tPV7pwSWmaMWx/IDNJpsCS7nH6m/53GSD0ZOkZCCL0A77yiBrvPggnPqQENiIzgfmIRuOfzeXeOf
GcoyxZaJ22AZGavDh+D30IRvBtFob/qfK1lmxBMPZnk1q5fbpx1gJsZFHKZ9g7aBsjn8RCRnx8TH
DiWjMSC3DGof2sDrbu3xAQ8eNH1Yh05hkuLrXS66b1tqBfkq4esy23qwZ6U/8h5WzniatbZldldW
AmnjP3t6vagBdoSx+AoDlTA/jOCANQmy0GJ6yh/+wMFC5SrmrsYuklUYdWgVERjGzxazEAcK7KKJ
KcUvId1s3wb+X4vpBENRAsCNjeiwNQmPRpYTe1LRnJqAT+57z3H+cOPkSFqlouga9AjE2UVL1+0W
6Y+kfxrPnfCukooSgpdmFdcKvLPnQA2A3dX90IDBRntHcJu8uMUQftzd64AsfCJDp+Ibi943PtoM
zJ8jLeoPas/chaHCcymrBgnzLiN1S1HvmCGaL0SGb7RIpFhli8ZH7t2oanZwNEGWJZSbFWKlWjSX
b+xjSg88aZjk2wOFi9HltKj/OP/qn4TVigFd7+I+qt1aJrWFURjEjp2nk/tDVmC2yshIh6T59n+l
6lg7KDs2jqdMl0ml7sx1SKFlONzV67tAEsxIvu3GxQVOePudLDmEXiHvffhY1EL0gbVzf7jbgei8
uVvygO18myikGKlQSwQck2R94GD3XouFjYwtvVn1/u/3QhIASJ8GVuNQ3kLf9Io/g/iHZ0x6B4MY
mLR/vwRcr5hjANerKYaSrWBBFZxxuNJPJhpDgxlbR72uzaT4ES+QOrMViTpQTHhRx6Dy4m/y1F7I
DS7qlhNrywYCQeBjn5RLvTJ3UnwqpLNpV2lR1gkaIQFMEnxalIKrn8DUdR4aSt1R2WMQl+6YOaMV
2dWnQNF3B1zuWd7bllaOv3kyFB0TY3h9H1E2jdb7/DOad8ytFv8fOWGxSheJ0D50L/Bm2VUvTyb/
jK7P241wmZ2LzHRGqOpRaWsfR+3XTLqn5dffOEI7Zz8VrIA7/vKg/A9dUwzbA4CkY7x5WiT08RyM
Ap8ZW0Vy+fkanX8fSATqp/s7AKs8+Vj4pp4QKyaYOJqAkT64MNteuI0fL2gLdHbdF+4DLyV34Izw
pPYDuTqoiZkVOojUBR077+3hjffkedlVZMzjKG5xEY3HMBv8pCqQqHY3gaJDY65dWuUBgJ33bLV4
UxHhwk1kdGguCCRWBq84IZ4w/niqEESO4Mlw/bG4z9KnLXrIvaA09rVrpe0+TynGwx9IQDytALR1
hMgiPaWnUHo+0DnjTTii2nLyvNDaUp/4tCj62WvmHUgPw8Jr8MiXVyFaV0pzkhOE2BkSp2uGLMSD
CHxnHic+glEWJ6W59hzUkpjTSTu6BDC4W8BX5rfbVVjDNfBZl0ZmQ0fwCTnZKYoBi2ZwQZk83Ddn
ROwr6zV9GPIosB4Udscg/lqtf4EmYFk/PIA3C4GoSuailwIFW3ISLhp0cXDkdf3n17wyTWjnwlY7
v2OJeIkGkiGoAJOQT919Gfg8bSp5jMo0gd7C3oohbjHUnBAfewvslnWLx2QmQTG6h7gnhiw8xUpK
Lh66yA5PCHQmdi5CJBUUx3Ol1SEqE6YcgeDpPBHD3BVE+EDm6Hrh6oTkd/0cvGXj40QCBIjBn4XS
TTpVVnRCQiH0AhuDqvONLOBwOc1jqJmATLhD9yKykxP4wKNEGt3Nzcb8eQujkEArby+cc2UD6FVj
h6EFOCJuh3N+xgHh1KwacyxzWJk5wG5M3WNRvGgqKfKKzKXBRmnV34VJQcVg4oJHZIO7TipZg3dJ
YdkaohEcg1gDU7LYLYtBWVt6XKxp0VMajhCWfUmQUG/xs84Va6rxCKpJ3Glm6vLg187BvyoE0Dlx
9iHJ2+5Y/oj66AwTLBh7njKuzDgv1kAIcb/J0pnzD/a5zx7zeLp7APxtlzIiV2CQqGvKQiX0V122
MH2qrlHZ1E6oAr/4mu+65DyAO/nwqCiGTClREiESPZYI47EVmQ7ip0kccujGfwdYLZ9nZhPH5GbS
sWpBy/c+KmBTh+Y49cvrtrVvOtG386rLMyxeb+vcGltdc4yhaZFA7F7xdQgP/t7i9QrKJgU58Bpr
p6Kw51cLuwrmp2kLK06sRnuKhNCr+2JZcQc+kSXb/YwKG38GJ73sAm3HfKlO3MAzxrV/xEJqTpSx
/gUhlKJfJ/ZpKPfW55CQWtWIBT1U8QxQA7nuY0E90dE+2ahpTnTjkU8AjaDr/SH7gKHYjs05iiKg
LXFgJW7SkPTfpiM5ltM7ZPSGjjArIbk1HlX88RpXUlgYKWrZSKoNOA3OMuC/w5x0LxTsScx9xZQw
30pND0b2PsV0z1At851hnNE7zHNjjO1euZ92EAXetEJuRtMtEs9gl5EaoE3z/BQ7uAmjXOLWoAtb
IrcShp2WWrQRCPhM+PYyrKmARP0ROO979vlNRoHMNOlDKopV/N1NPtlr+vLhNMcaFXWSct4ICa6i
r9PahLvlvxBI5E0RiyvNbKx1pZbnmkGGuO2YyJpTe0W1/f+jegSjkUQn8QfrJNeuAxVUnsCprtu4
1WcbgOqsMy8G3oiKilHG1EFvVySLAJcqXK/ZMaH9tpIQrJmrtZKv8gW8o9/YeRLLHGT4iYgoFlmi
gjJwGnAvpPUN+g2Ys2ampa9vz0Az/Kw+tzSLMFvU9g/odOz/tFratg04njommAs9M4YuiUsN+Or0
bUrjywiQzn176eBDR3bK1f8qaaO6Nm8hb3R59zk8/nk8bVca/RTX0ZKRUeYjXKr3jxRt/as2oLEY
emvztgfaOPRZLl1WfpLAunYm67Msh0xTOP31D8Zy9uFikqcpqKmVU66QVcb51xbdf5r1ivrZL1ry
Rfrdq+qC7Asw9GCXwfupIORnHYyJI9r0GCGgyj74HhdIc28KzZYTSFnWRn9gGZpYdwHg11lxJ2Pi
b9xpZHU6q4kqZVGojxiLFmVjESez4uC/91yQsXdh+9ad1Be0WAyQULrZTOBmrep1GC/qE5oBf7vt
z5DrkvXBv9MOpCL9fMPB0mk/uf5hzzJJjYk0SottC3xL8AFPnevIqPZ4IlUm+g9iF9CIOg4vl0q2
LyzOybOJmabumtcKxhLpKm8dDSVtazCBYocyx9Z3S8339CbG+3JdT+nUvgn5Uv+xOjEZ761cpOJ9
w+5cE9b32nQVisApLrFN1pH2Rqlj6INlyM6PyH4bYe9GJwJoazxAkSYJ/rmYMEdOLePzsyaePOax
QiQ0qSevF4IpFUP+E3M4f6pDCp7za7yd02MHQQTVmE2yPLFXploNBmdYkSHEK3NieesWBOI1yJYn
vWbI7LNAvDpkhrFrtIrYUXWmG/18kw1c7/B1rVhyJLs06gaOPARYweWfkwnzGdZU4ortEubBpAbJ
DmiD2csWS3QL+CmfOS0fscyxcVmKXbzPFE6fTRvrNm5DXtKG7t0yXOXVldZycSS7WVkJ1S4qwDov
Az8gTRoCy7NSykzelnbgSb4x9hrdDWDF1mWu62cdtCXPLVh/khJrQ5aQglC6mYv72OKnBa1QU2sP
TYLMlvdtxuDy2qwArUDiy58lAM4yLpLZuwaHdh+Jn1mb309jMb9guzbfTeT47SY2XosLHxrRlfxR
TteDRPn73AfcZT49eJ0Vd8TQGjbp6bjEFrhkpOe5ye1VQKljxAcONLTzDC9KzyFeOcATM0norRSo
9kdvn5NQYQ7kfYnGTJgy2fBAXIX38izwYTW9m8cCZQtvnZl7Pt+03ggIuz7OGV4/M0NP+3VVj4KD
rgYl8vFxds/cA0iTiG/6ve/J7JPPD+LffAlgYHUefO8gT8yI/foQ0UoWch6F27kAZm9lAlz+8+nL
1rxBjKI5+/6PFWUkVAtFu2Cs8AWHWhN6Ta6c5oOlUBT4cS/35ba6OqL1v8kIEFxggZr8D8FkOhbd
WxWNmvjZy8CZ9YgWMS5p9P2Z3kvNCvKT95o+edsrrVnjVinwysC0jLkYrenMFB7xZ9WttQqw2Ji8
jqzKUXtGVhzG38v2YLUMtYhO8apK964sfbrLsk9UEYsRFjGROjm944PfuhqDMoR5MRCA9Vpbpj+N
mWe3yjXVQbeOSLjx1FTkvUP0aDFAB81zCy27zgkoEg31Jupct+fcAqzhSOOKoAQgaAVSIiZ7PGNJ
TZtfpeeO31U5H6RUQ4BBbFWNKB3myhcwxj3vf+wIo+BjiKMTVjb06+NMLZjTe6msoR4TWBwoFH0n
Hgv/hPS6zAHHY69sW+AZFdaac5LS06KN0WYvxQjVakyJTRnecsCbDpQDoBfzw9xrpTJHUKd29nPd
yHHoYmNtmDZYW4Kn3eRB/jYo534drB7s+g1yzF7zMZoYLIIuzygBsDYNHUsgcl8OCninFiTvYaQt
TDz2C3HSCHHeYh1HtiM7Utb/lh/1Tmp4aTaV79XclM430g/KtNtTvqNMkXlEWNyvjcF/iXjSAfNa
smW7Kmvu1KduqsngM4icGkyPs0EmR56Es8O4FkPAC/m0uatRcRBccFcRHzoaaudfWDXJ5TZDAVq3
DqVbUcEBF6iPm8rTvXq0P+6cXvQZBlcb2W2+wbamUBEK35y1V15cUeb5KZYzKuETof/N2XgjA20C
Yydtrkx5gGFcGe1DksszG/IxjbqGuGr1MA8P+o084c9D4vr5peVyst/ImiX4YO6Fq5AbNPy1BFOB
1EAsZCRk2jIk+JZ6oUtdfEb0WDSWK1BfTblaATIPlNK/1D4jx/CC6hn6f/BNLukC6Sd4VRAlHU7C
ESTun7XRi0Gn2QES9Z4nTeS8BzuNB/DNhr7IwxxsV9Ps+B7gGH5KURzOtODzQ4v6CFovxiYKJoxS
CokXuqxp0CmewmsybltAQSnAoMHupLG8RuSr1evqS+Pse6tCP25Lxz0oM9OwRnb37SN8tkARCWdl
jxi/C7HZF+XIKm5HKMcgACOe7OnWJG/qJ07mn76m43gFls7xYSf+dgE5DXWOLbbjkEBObrK+2hiN
PpC9rWNKa3ESxIB9u+zMwlTTNa/99RgotF7ObUmntv7ChnTEeNYz7RXxtSkZQSjvOgPcJH57uLPf
2llwoj4MdLtBp9BDYuPzKXbMoNax4xW9BDUrd1UqqcNZvgUZ5xqGogtx4J691z7/omPF/C9vRs1K
WusLNsT6OFDvnL34EO1s3TbuOHvbbF+ml+PQ1fJ3S3PArF4gTmQCiRmj7Y81Xhs2D8JwRTfdxWPD
GhI3gapJljIT14pvfdOStGkbzXXs6sNeeHMLLGkzYERLOjzWePIXOpi18hO9wncw9va2ijIor6uz
C7eMDhV9mbDofBCXrh1+ldn0LCF+8uTtS9RlLj1V+/aHhba+CAXc+zBq7c4A6flYosUx6PJhktVx
TSyTEpJ6+39uj8Ab/i3Vx9T84ad/ZBI6U8+e0q0dsXRMDW2xoHtkctaTgMpqbUNCmOLpXsO05BsM
AYyaz2jz1KBUefh0Bs7N6q96fLsu0QvS+YagpDCHlSvWMuZIX2ceCpXRsb6MSXftfm+TE4kaCTmB
vHSovK1BoqyxNR/NvEq41e7GGxsjkqxdKZZgbirxwRfCum3AFqBXqTIDdX5wi6edGzz6DD/Ozv4h
bKsWfjFueIDlK1JGjY9YTxpsoQwBHwORV2zWxllhdu+JS7yabOx0C9BX7SmbzWXcKUE64EgB3U9H
rYdB1qcYUksxOn+1OGB3diNOqGIuTazH4Hmm5SlHC+6Wba2vB4BIIGwV0KenMt5DtqPLB58qUjxI
9k2bl46x/pMB7/aSkdhBb8l7ih8CWgjKo8dJxxsTMTyNNVX5POe/mPh2TtV80CfrRths560ncLWt
kBnqZtpdjjgVf1mXa7LpJq3EDTeFfFCkCkFXoz7cG3QqiPvJ3d18h3AzpTFpqhcB/ViEwlsRTMoD
vyOgzDJUMhnp4TsRVwI2+L5WT0mbVT5WZttdhJ4SzneuiSshIeL3dANgkmLWD/N+oWs6Vw4iln0n
gxXa2sOkPErhj5SOGqmiBJlRlphChcPKstyvIHzBhEhVPO6duLfe1fx1rZ7Ph7jlE0hpXMUsS/FQ
Dv38pBg9wW0deVYE6iO1WSBlcfRw6u3vA3K0KCm87OL5IRO7SS5P0mH4YeqJOtPk2zfmDCZZ+NeM
ImWkiXmeSPmqdZhp2uHS3hT6G7+HBUArMDRv+PCxbua4vot7ldbo4mxk/jVZ6H5d/shvNThGWor5
EbCXhUY+8EKu6HiWFp2K364Eeln6ohmdDLcJuXJskE3AVa5/q/074fTqv8EqaCYlGVQcjitUSQSx
TQIGomn23xcYDFCmBFrD1uz8rZn6Wf+0WDi9mE+5WwHa12cqXkeCBINBvlXkwo+Y1EpJCRTu/N5r
wH6RIhWr+GSOTo9yhy7zb1PDG8Shsgpher/xkAxOVNd52Q6GU0k1EL4vVcUx0sJl5hF/fISWMIv1
xjxUIFaflZmpH+v6erqnn4JLSrLSogRDaUK4wh+VvnNDep4ZFT1nbHOa/bOnQrhmPMFexjLE6NxO
kSXw+a0TEtf+M8ssIe9z8+A4q9lYB0/KZ2ytAuxiNmlb67s1fmasa6WzWSeEcCyQ+AhhZMMnovIr
Ts1Od9JXQ3dLCojSwuDPXe/tkXHHfEEMLg84nso7fVkD5Bn3+OmdzhWk6b2llSaRW/jeOWo5QSJp
OVdVYHLJlpqoo+DeVFys2uScIWrRYDAU6OoAFyZEYZVyc5E7oy3+XdNEmKUo2tXtddRPBhX6bZPE
8YK3fVZoAjNf9D/PnOxRV5VnkOjdLkcswU7Za41Wkn4CDwX8LwXASXIEK4RRK1OEA+4QGkHixRqM
3gbTbI99F2QKG5Ubu5HHOK6HVcfzKfjCd2a0/PeOUYcx/uyIMYqFv+sIJ3VscUjnzItHV+JICYQT
98X0bTlp657pTVwZ3uugTQOZmtDztvtasCKXIWw6XLw0qbJ9fUdJMpLIfddB4ZsbP2HaIm5lULae
rgIQME8zoicKcyOa7URiZ6kwtGcrBD0dEXL5DUF0WU43Tn6ZAayqFl4HdHHQZcouBXsQGoplyyJJ
GIFU6IbTQyjCZww67mlJJZI55lGa+YMkzaSjhMTLB7a1tQ4GRtB6cXgz06uaHHdxCSOUwfi+KLJ/
GxgfDjREwk6Kzzajx4xBioZs+pUa7EjNLbNCy+VdOAOr1g1ls/b9C9mBNmsGXrs359id8+C2Kr5S
a1c1H76stTdHs5a07cYzSEYRHHNEIEFQPN4CZ9qIGIitMxUZQz0bXDij+EQeZfs/mVKyP/+Jrfn9
5le9JFlvLFST19zR5YRtkVH4VKoJqklOXM0q4AhW0usYNUX/kaNerIeYNhzeatKnsA8o1zACoCqW
Jdza5TNVnvbA1ty0qbS5XwYt5dZejTQuz1mdA4l2dIfEUT8K0weFqrttPcpEgeU3HQn0RO3lYUXU
rpoQVW01ydY+1/yVhB206XK1QZy5+M65R1qkN/k3bIWOM5xB5WKNE10K2bhlbsAPhF2ZmnvZv8/a
KQ3sio9fvu/n1DmGNB0xwamH3qLv8FObbVlLO+J6ObZQlueMFM6vKfr1TrtUMaSCWDQmlCVb1Kd9
VH+dvU+L2J/bpPRk2DTAiC8EhVCKVLuVU6X/qJPdaMcdNUK02YWYg/PT8/ZwOItNeJElc/ealnol
UFikL9DneXWQTYoMMLB2gUmoXgtu7Pt5wUifdbC9s44oPanB3zddUMicRCcpHNq4/DQFZqzl/xGV
rEiDpCa2z1LomsWdwlqoBaS/YIjTTDXKhQFajVTQSLHmDTl60vepIwhpaGFDstLCTmdQz275iTGB
DVR77EJ0q+ortb+KLvvqXcGqhRg00tcmT0X9AXbDBCp8iRfCyJPMjKO5ap/ZFDsK9oITMO4CkyI3
Vtsl8R1BQoiMHbkxZJpooIoAzoEwbadPTdnFPJYx/K9BfxVn8mb876Xxs/+V6jyyeU+TyXsEd+Kr
88xYZyfknaMYwtlibmeienvEeYHrlo/Z3B7Gwd/0a7YL7RxgC57a4BaeQTqPx7t0QwCZLkVeq467
HQXL8DMzYoVItO4LDyp4EbQv09D3GVyVRxGF74U9BJlIF0GEz8RXd+FvqaY3FoT8oDzAprW1qTk9
Jv/GQFKJNtt+YnJwdt0FXdgfvCilIKE0Smu5NU6+hiHWU6uwakioWbNyAZaitMGt8hrtABISfdQW
wzfSYnVW1rid2rtwyGJdJIg7hn0HaqARtyg2avYukZobHYNPEycgW+Bzl2bzP+ateVBNh/VAaJ7P
ySjxzTf/AmXxKxQWMZogxbWFy0LlJKpStrzL2D16criyxH1x83kudkVDtin1xSNwjd1QYNZ9Ci4G
o7f9EeSlR+4aZEJfJTHPGie53bYTO93vmc5mtF2ohw5f6Hz/ucahixCVn37ttqVXIYecnkwRpQe2
zlzozuVpo68GAIe70XS467eBB1L4pwcryKpbU55o/bdyFbNsOrXimhg6lnUq1ChjGXHSSgLX22GH
6urvPqSxhST6ibidEm89tp1CMz0l+1JtVyBisj1ABOtpNjqAB4IgS43RH/v3+C+oEqrnka8GHuVx
QhXlnL//1PjS7k15mh1b1MDGNfrxVyFgvTrxa8Mt/R/QpFMXDod8+AnhCNWFElJO1lX+h9f4z+te
+/O6DBJXR151xO3a2FODapTS9h4Nb1xslLACYfPtwdty6OqIPQjgDIHFiRoz5mErWB4s7cBdKXaw
8Tl/u4GqR/k5bvguv+lcSqiLqcdbzomay2c5zodxUdNEKie0BZAoenrQhH56N0c1u+OkBKgr6QYM
zFZ1X8YlIwf42QZ0rZmCcmwFkioWPdy+pewGDswRHG+6/thxHeA2x99mb1ANLVubw+jvPvUvaEci
iLkyCRQ5LnEryE5RnwrzpnU6AKLyB6UcES3/fTxgyDU1/ev0MXplzI5dGlUQHtu97SOe8Lig61Vw
SQB36K76BFEG8TdFphc4i0r8X/plpdid+FtnxUzynyWkIvMEck6Q/WctyTG+3Ah8E0acEha9eR2E
Xi6A8kiu+CRogiTZBmgkqAe2BD5BuoQGp4rm7DurE7hCe3MtylBeyuGtzPYd4asGgyVME9WI3O6A
Ja6qdCc2bTP/Rnx+TeO5NSyDIgif0LBsHy9fUm6Xbrkv1ymqloxJdZbM8HdpXJa98Igi9jAtyiPj
rJ5TBm1rtKAmCXrdiEk7UH0HRoBkThjAbB+XAgUcqVrUFy/hn0UtBCRtEfujXIetHv/AY3JI0dCb
4RiyAa3WDZ+30QUTZTxSw+5N28cLHgwe7ZPkxKGZKm98y3u6AzvovaDaYjVbHppMe3OxDlr2VTH6
zg+S5QdZkxFGRuJingb3iGfWtVbmHz18pMH8kpcvw3IINwXJqNpQ+w0GBRrDErq+DOomU5CBSap4
zcy9e3wbPrkK45p0/vg4TDFuP9MjcCaK1kpm6WSoeTxEqNOt9uvuRHipGNu5q9TgZC+ShaUcn4i9
szQ2UGvHQK/5OM8ivkMO2loF+HZFvUzvJXnPM8ChGkCdeZvrEhqxdsNwdAM2DSOqFnG55SzD/JNc
0jvs/Y7tTod307OHM00vGhQacujYQZSYriHVabIXQH+NSE0A7rRD7teOqFbq0Y6UwjEA2+hPgjgM
MISHseQFlSc1ERdL/0+zcGGLz0aWA7/cFddyzZjez9B9Q8wrsdec7JTCdaht7S5/qNCJuMA+fSpG
SehitBD17CCW4l4r+Bd8wWokDv20Qn5OJURUXcvw59WBJL5HrrfjJHwRyitf0insyl58t+TrPqeJ
wXFifsLXoXG4yJn4rKhWf0OND5uAEc2yZbaqa6fnSCy9X+91JuwhX65Ldrr0j8smyKIsANjiGhe0
EoQk9URfsZ+yLguQIwJX/ZH/AtKy0S63NBLo6t7UHHU3MLvOXp5mENFXxU7JV2oSsMGLGMj7t6it
qe+T1RAeip3fbzOceydguiYyc0DF5Zq780FRuXg81KdS4wmth9DXS4BFWSTTHlKthFub6czFvih2
FmxjP1R4jj3KcGinJ/SYcZCTb+6b8Z/F+atw9aZlQK3sfhZkB2p3OjlTX+CTADurVjHnMWSkMGY1
TUDU2mBgaViVJIwusOzVpwq0luRJZjhzEFAMBMs6bojepH77drBjRh/Uf5w4E+hZZ561JHtTSFxv
QQg9hyxG30dGZXbCL0T23fdQnbmUXu7iqcyDg5x7GUcLTxSW8r3QxdX2EqABZDYM6pnBf6qQfBYN
+FECidQOx1djcQGJ8tckRnTi4IFrIU6Y/NvRfBOubw3nvJNxDQav8hRxkdofKBkZL7KBGans7PRa
BhYqcmqUANx8CN7wbricBIZeD1E2/WOaP8Okx81z3jM4ybS90/2dRt5AAAUQX+V/tS+1h7l0KnKT
98qSEwxBeGfuDP4qDR9t9r4CYjCZpuc0reXezbeSEboJ7NfKCZnLNVEi+KQz1DTbCOlCrqAFc0uT
gsZVFv1iFuKugEKrS1HWJGH8mO7vepAmuYQKLfDi+q5L4r4zf8jxxf49OmGNvb8athUpSdWJgs10
nrqisjRHmr2rrLHI9gpmpRTlPcLDV64rLIdCw8zsnnLy6NvF3AMrgmAjz0+rhXkl95sCRWszgUT6
jPhrZj/VJLyeev+EQV+AUIh7i7GrHrLqIUpvS0HZWHyEYXZttimTCHgmT/lOIefIA9W5s8ffIm+P
Rf6pDy6NDTwkxFf7gpiGdpIy69CA7d/dmLywvMAt87ZHi0QOT3iohtgiewuD3iLseDAExHUNfHAU
SrchJWnjWN6zeOgyntEES1BtJIIEyL1UkbyxRbx5Ciinb5zS4si9Ao0AB7+Y9SezaiiBSrxkrpm6
pjgxYxtn0x6wvjIjqEicgmO1GKjfScNg54/eCPAZN0C7EGUjfRpGOpUxxdsIpNVtLcUp9UzMKMma
kDTvLN6oqYG0J+SVj8lI8TbZliCgas5AuPnX88IhH597S3HRvp5p/96DNMXP23JgdlP2L9rOVsyL
wpCRr1bCcjADTD7aUSw6GX4ddz1ZaAS+iP9s91qDSrZgr9DPCRKuRya6ZAcC3x3ouFDsOkj5xCHo
PayWX9Zyd+OFkKr0HtSxRnPuMseNIQegPJgNC41UJE5o1oloA7PsGczBNJtcqYRUHJei7PBRbOPP
hQqutr6LjuDtS9dXqvz+kRIYRbjg9o3cixlnIYqvYPDxA5tlXRvQVeZsFjzRVGTQ9o0cFjb9J58b
s6rwoLBI8X6UWiChb+d9mTdD39GljyJs5xxxtZZbolxG1nRr1y48tRsGcPQMTxG6upOp+EMOCxDD
gWgm1pZcjTgaEQo3B7l/2TJGXvstcv/ay8m8Slilo/6plPjSs+tfeUVKXDSrXAwYLfil2QmPUnt+
Entgj/h7Z/GvqbQxRpfKKneovWb7bE2cxJdIruFzF/UphKbnVc4Yool5xQKKZw6OvDwTCif3HggH
KzjfG3Bkbm45SpLL0sBeJMhkuOtGjF6677I8WkhRzuK+Y5C4QR1fTUkJ7rDIVJTst7JSCnng/dZZ
lz+4Fd9vbJzcYpIKg3Or29ixXG8Q92sj/fwdb7BWIEA9kAJq2r+3eTmp2lJTElUIx/S2AWN9OhTt
YQcyLkp1Yh/wZmXO3xGp8wz3G1m4gW94Q+2ccBhm/qJfBBTwoRYSWqLk+U3FVGpbejAHDQc6H7OJ
iWArbZ4BB/CNiAC6Lvbe3jC1eL5JdQa29q+k6ru0pQVmlzUrNK1b9l935KBImsuIVhcSSVMd7I0A
d/jKlF7Q2MAOIQ5QRPNG1VXNEJalnpwLXUBKTtUqg7WgoQdod6ztLIgT4oABW/kKsJtkLDfGef/z
1+T7hl89q99+HE67a/h2n4JlR+Ek2FiIas2AmMZJgZRvvSed668Y1TTkG6aElx2TdukUDIMIDX68
847Aj6xamgOZFArt3swrSsHmOxhSBnCPl9dVM3VvEBT+Rv/nRgxXO4W4lxTsdNWTdnjqme4oGyT9
RtwiTzMDDa5Xdl32VFV0NfXP1dXrK9kcyzkalidyfEbSZMG9/on6tuVJbPc4qbXtBojhbkwSMJ1x
OJQPnTps6jEYsh1iIs1m8LelyM73HMl15RPbijthnMVeAfv7hZad1uyZcFCPGV55P7OWzlMAHGgy
LdAo0TuVk0YyfgbRFAKuUMSWg+8DkcO1TKrGh7iT7LvaUrRpbJprEApVwTq0USOoFGyxdX0p7VY1
J7BQII9w+wmn4FTCSSuBW80e5NFPk+jCeaGyGUIkb5B7KllbB7Iw10CHpaP6VZYYbuteZpRsO5vn
PlCWOGQKdH9WCI3a8DMPxTV3MXIV0bK31aK3KZsE7trTQhA371zJKeqvn+Th9Ab7ciiuEx65S29J
RYae2mOYTJw3U7CVRfNZsFOeeeIPSiWEuiN6ALOQb4MX1wU/d0AT8XSPjMhynaKzem+ByID8cMOI
f4i2M7gEzYOe9VO0xApgV1dDV+LKFTM4YkWHuN8PnYHXl49bzjL0S3z/IavnWluL3cvOXTKiRvA2
uUMsL0lC/R4i0s4xWq5qXuWuJzH1F884svg2xV6MxQtZxRg7iTgHNbFpJ/GBCVadsd/2vRfNdtX0
NQsGjQF/ujcu43kaQNX+0Qq/hBy5sitq1MxOVhHdqdgfzIfSjTnm9W/8S3T/zaGiSFd/LzBWY5KT
cmV0tWccmdBNGJfAOmPoXsWqZtx8dUfIBIm4Cc2ZFW3n4j0zsRV299BYBuG6ukztYLC49Bs1WrO9
mJg1v+XNIfFY3qwxlEcp+fUB22+R5N5vCa0NKqcG5f55yiwAY1GwAmvVeLD25SNmESTLxNBEtb9b
LBtDJu6R9yfybcs0fN3UYP9zRS3xlJrOYUrGWbpET+VTZPWRAdmHJ3kZ8WB62CYf1Oc5cDToCuLl
OmLy06ZoI8CnxOjXS4xBwJpyWkK4yL/Z2icoqviV/JrBbvnk0wUayHr7KpATL32mc+fQGWwvU7Dd
wKganrzFMZnMxX13FLWsnAv5tP5JTW3vxyaYgTHcPy4xpeSFdBiN9WrmndX3+ASY9m4py2SDCHG3
R7YB/Jr19JMFpmMAvBwAXzv9MFFCZARP222c69yPLG4lzmspFh4mHiwPFC6FY3VeZ4w+SYl3OOTB
H7mMT3hRt4bQRSKL5OyiWP3D96fI1OaSJP90xcqhZE8q+8Kpwg1vKcRDOv3aJqq2maJSn71WWQYW
515XRLE9uMFN3QathgOXyWun1ZLL530Ix6vey8bDdEOyinhS+Q19GTrhfYreF7iyeSjhy29n8k8S
q69zqmUEVQQjCx1WAerZ7mkOwy4tLebP1/WVqXPZ4QcrcFHKzeqCc3BVq+Sg2YV/PtQi1znK9gbT
3yoN+1ZCCsd9fpm7gy5vpDI826Zehwvw4aR0s0lOjHQtH30SSPVP+EcRcR8yeGLSmDQzYm8etn03
xvldcFyBOfu9on6cPwRqtpSwMfvXoEZvrjAvMkmSwnMqTtOlGw59MaFImH0h1zrBrhibQPduI6eH
u6kUxhfTIkSGxbOX/Roxp+cFfvtNekIniC0T4uxdvl7/a0QoSu/5j4rQs5PyMNzGzlzel7U1629c
b0GklSVhYrlvmikwqpRz40nQqkJqTn4ZIEJhtpo9AxAnEE8izGhRZjzwKWV+8VhGdk913tZquvJP
OAefqbCqQ9RM02sLJOTolJg9SXAOtviLG7Py/gut0NnT8qdPxsxZPBQA5/7la4HesDCLPuUcxm/h
9SdqiS+cilo4U5E9D/Ionn156B7dj/JxrrtEX9VnrXDwiwWOd+foNz6ApT2owTHpII+0yim2cGKF
gw8L8xZZSsnZ+gkGZGfk2PS2VQdrq4pkieqZJewflEleKAjjzoFSS8yQy9FixSmUNu27oK3Ere4i
3yBCPKCCyOc+atniOwC1mNfjmd4mITCtj+cPBcrn2SOuN2S/rJKr8RBCyrotWykarEJyIv/POUf1
t7YW+2seP2XBv5CY4sKd5VKGpKRCdhXJMJsSJVgGB8xL/VbIYkAA04SjB0RiY9LXZJTIZqypXM9k
2Ce4v/LxJYTj+Y6VAOUwgVaOy3R0saJfKeJ62ZB47690z4e7wphT3V0ksiVEq3ZsCwVkrJ/Hbi/9
5wfGG2KQHf0SQzj53tJiIu3NRTedNH5a90UQS8SjISl8F/WPXxx8W4iyg5T0SQ61xLMhf1R5gohb
EvLj1B5wfCoVTQkt4enoNGHdNMRbnjGPKPnZHTvCDPFQTikV1BH9oU2hkf8DLoCdRagzathHm/PJ
Ps9cnjFCSDsI1S3lBQLV7lAPYoeYAZIkbVumqRhqD1ahiFNBfD5mktONB+q5BDAPHXtnZMoz39Wx
u52lttO9rfzsjMxVU6S3nRwdacVMiDujYzTLkJrwpCzfQzfxy8LG/Cluz1VK5ADikQn/7H3KYTOf
J1gw1om7fbD1KPWuX65JawXrOicK1EOTjkb6hqGkkVeTTSdfXGYePDWcM8BXJQSB1BEbAbUA+D73
3Q+EXfPe/fDcYLeEkdV6VmyP5MokHIlRzEfhiHfAblSzWevF/FiZwdCDAwRj8a99JZpfXuvIvDJ5
fG1xAjrK/UZxVOuRl7p92nHlMZKlX+AxFO+snxGqKpHLre7sMk6Hch2dA2cYv4YTREv8gm0HZ9JZ
k4EII7wLxnD4SmIQ7MHY5aDGfj1us7Vdl+Svzxr3mXZ2ENwqu7NYW8ixpoe9j77InvV35JDLuRCJ
Va+CMOX72lwsnZx3t3NWrSowe7G5sedpsqA01w97shAPb4VwH8L7Zod6cOpF+kcHf5Bv8Wshlk4c
GteY9o1zSohWvBYOmDmPao8r1dcke7WzUcOzrk/7hyWzCDqQAMYI1yMi18d+eM8C0o3ye/CKxgvm
FHGtpy6m9kK/f6KxgBO3WLu7DIkXM8poPH8/+aAyvRQMV1mqFSYpRUCHbXjZ59I+4dOX+pzJ7SbF
Z+M2ssRIR/m+GbxT/XJRFUUaH/QJsqWDNLe3J6eutGOuajEXWTDIhvrpp1YfbaM+5AjqNXBAfrBq
ZUZxwTxNT17rj2zWmcXBwS81ttvE4StJrQ4Upsy2yMQB/6LNtRzxyxJjuxbSKxOy1NjYgujXenz3
tgJL/EtIHNHgUcCsQRj62QIjMT6mg9jEvFpgJ8Uxetai+9Rndt/WBqUKg/UQ9MegJxf+QvwVVE4y
qU3fS0vOj4Jlciybnqak03vTSgDkXs4vFm5olotvc9jeqqKAvveTkXJtQtmMhtvEFx41Xbc38Au8
2jC2cAYblPrxiA8y/dodB1qpRBGNRNjlDeq314sB6TJPxSq8H5vJwUFoykbb4rIxXsHYgWnQMLEi
5bP9zNrUcuIBaBH8bT/ZQr7FkuX7pBpSAXJJGNr0GlwuxLbCAtv/9Ih3ICBMzqJzdj7ozDCEYA3Q
9Zic9mtQveUc22HJPK7L+CZwi9BO68z5wpdljznPeoEzT72XiiBPefkWUZW0YmQbqHSrf4iULeLi
g4l1tMe7W4eNuGQFSWB6P9DYhiFtMMybf1iRKngUrNza0HGyIT0y/cAUrAbeUCOrYxiMp0rW9V6b
dApsbqmYVMfCWz7IsjIPFEOSTYehlfFVCu29MqSgydkTHV7KAepyHKSp+dSmRi9uKLsFGGatMYXh
dAPih9is3Tx/HQeZWrd6SpXD4oZPeeL9zwJZWQlKdrrWvoZpmWnTUEBiwXBrmZ0L6O3cwLkeJm7q
fvA/rDLJpJpmb4ldX+iF8efaUDmYq8f2D5Ay6UlXBMO3D1tg2dNLvgApEUdJ6zBjtiBCuUMAbh5x
TAWPk/00ihaeGMLaTPIE8r71R6IQBtV5ePNhGTHM7fvQbTmLJrF8HCXIH+XrTwxBALEaFBcK2ziW
ygcjPcO4ADJBTp90Hsh0csTSerOdUwJpCtHKyRiRB4p+3cMDVy6icnQ4FddwgMxmCE6YesNSWdma
tbYp2Iy4SesAnyDq75iEvkfF5yn6WG117xbvhTQ40KlKLHizDCzGz8y8uDz5OXGk6ZuGuwqM28qe
KjhIJVFAHjZKhppd3GxCDy/4RB6GDlerqWXSujYeZe49/LmmXb/v1TrJ4uY0SgHC+cIuvHZVgcZK
Mv6zNT9uBh273iNL6+nm0GRfpOLIeubUqa8SECZx0F9YqiRB4VVYrO+O9uGcRmA7DF/iv6o7GatL
L+F3jxwtAPtqrpAk8cVsQ7MCKwRXkOzHzf0BA+NP9LoSfTUjszpfCT9m5zuKs7haWHivLvpOMG5v
VMAjXhQCSf/Nb9eAiS4Q3rBxqLA7Ce8TSTrX0ViCvXSnwgz8s7Vc9JsB0U9afpG2Y/6pp4KP/uJI
A7MfThHzs8PDw764hhrIpMDpw+nsOceLL8dBjJjIg744fKeSnJ7vQbOaw4E7tXjYX5oV2Coh/4R+
HTk5tag6dQTeuPfJUVPaS6lq6Fyz0vCO/DB6vKVXqHuUZe7zVGTRCvomqt+ud6h+0W6hy1pbeFgz
ydF3sX2FpSZ6L79jQvtJOnhvNkqUDw+GMvsulv5bBYNaTP6awFuz4kcsXOf4J0oUxeDBm8Y1to0E
GQXAq6IPE3hKm8y8POZB6BSfOlns3vXsjveVLiMTTiWT6HequObFePneahc+axQNW31I3g4CPHNu
mw83+sbBGtUZOyg/Ya8pmfv58yG4yWiD4/5BbD2CzZA/xapuuU0EaS4Y4gGGZA0+qlvR+YzoZOpQ
hJWtvqvhc+YuxqTJ16w5KY7pqVBw2T2La5Zpoq5YmdvA5rvP09jz9DJsyrltS/ZylejqyxDCIk0M
dkSZS75M3msLgc2gIdPNGKSm0VfsRn1B6so/OA6e7ST+xf5WSOdR39fwdtCCUkbd8YULaTCS3W8U
QVqmPkPmInp9HSVSuKb1IX4rk/nDvI0Jxt+KoJqYodV7EmDYrrp0K9mbyYHSuy6M5apoYGWerxV8
iBZFUIXDHWPeUReMVjtnCq+EodpTZKl9x4I6ykHFfZb+rqiQnRNKYcC3y9r96uxJbNyaF5GNyv2R
FJjCbZRIj1fX4eZZ9cWlzngOg8UVF9pbmGnxne+WuwJuDnIf2fHxYP3KsdwpgMSsAaXl4XmgEHrv
gfPZkyBuKuti/ZVCo79Cv+7lt90U+zGL/gpxv+lXR5lKT8+XplKHF4x5vvbrWYzh+Ygd05gOjw8L
IUQOUK1EQAxX5NRWJTy2j1ZRT25eJIFDb5ok7KQdPrUVM730V3Swr21aHfw7agMObJK+Zwd5r8C6
/Me+L3TsGnnEhlLu+DO++XEloRpq6Fg74s85/5Px/n5cmneWUKIae7wL0W36znX7DYkAPt447YFE
s1XMeIZLzCQaH31Gltam4ovr9BCrKyOAA9Q0HZIuSLAOzapKhNYPyom0ZocV6AMLIGjFpyPp5fic
h5+dweMSWduMy6pOjAB6LKcCH4aI4FrU090cXb5nJb3DlA8xeoJ7sX/hFv7v7ekkcUDxctf82fVa
NzjA8a5odHzQEfJNg/WW9HuBXeQFTfnuicYmrjrKjVT7gA3qlqwqm/MRhZv2YsN/CyaNaDVmcwwx
WOPavrb5VvwiHGSu39Ij8cWWypwfFZhqJ8o3KB1rhBWmyGeQUiDa/IeSHbJWIw3EkItk1jh+bqqi
o6KWuHtCh1IH3bL2mnIgm6Z9jKNEmYHVsaNEjXEXbrwTddUUwrkYaYrFY/HvwrLecXN/6fKLpNpf
pM9ebbMi5jftXgm8UTHRWHvLZHeS/SViMK3CZfpSLTmVUbA8e9WIaZHnI9x+mgROkfUfAdHXlj2w
XsnADO4CWTLgK83cY8TFGTf+8cE1a6fPZThR5XU0OT4PlNl2HsrXASiZNnNnhL4bTkzZMRygY/nP
UAneLrHzXfRXRDW7V3Vg5wb3ZeISKF2Nqe0oksCTWh2gBmpSfQMVV6y/WzO8wjvVEL/7A8TDayUJ
HBqjEJhIh3ISujdzxQkqPnuwW4LHJSBIW55Y/IUTLSMXWNDIZBTT2ZC26L5Ygq4Q16Kryil+4CYz
Tr9fFvlJ0Ts3QS7ao6eNBP7KRmtlvauEK+5lwe3WONyrrNRV2AvQwbQOA9o1JJGss4w4yCsBftAu
4K4j/ZxqrdLSUigoIABP6oj5hr3lgz7q5+dylX4uHKkI2ALGsXPN3Lp142Cy/RwPY70IRZAaRsCN
LO4rtgIPzzvel6NvxIkLwPOzcItSCm8tJpy7IYGKQVWmFGpgIvFwn6mxfGJThZiauw/KuLh4BEvk
vfz1GR7BQHSmc8AfcA9jKyBp9xtiiG8g3JJOKVHcOoqY0DQPzx8FBWgabhyTO5gPnGHy9jhxWBKv
wz8CS1hGTk15CNQOqm54T4vaatrk5Q6qBB6R3zRsXdGJOU9aDZihCgERJmqKiAmjQIEXyaFsGRbo
RIjB+UEdJ3+n6/b8PLuvXVL2tTBJJOWyy4eGfVGcmAOXy5s41BxPzJJtZ4jkY15oGHHwMzd18UKx
WHhY+5r1dAJJgUfI1BaJ+G86gcOWOXTC8Nyh1E7cfdpV5gD9b2oo48v9IFWTvNx+XZhE2BuFs7uD
cVdSkU+V96nHI9wWtriDwFAuDrTEyHxSvyi3VF+8mZwO5RUkQ65OMNjTg34UAkiKla+y7wShDOME
7CvDOIjaMtuyEtCzmMa9fg61Y9mjmwrHOtybL3ptdWlMd5IyaDTdtjsRQRR66/nqcWqhlHledc1X
nOpbzy5MrrNxLo2TIKqqtHi5tnLftHrlHY+QKYa8DM1LO1+plsnuJbI0b4qNay32YhvlX/QFnVz1
WJh2ZKniG+bgMj9H2A9/yieWTg2DfE1ZM3YEXWP9Ig2Ri4N8n8bb3NoY9+XR0IObbjRGzvW3L5P1
dQ2y3rcTj9efpHFnu3qbUFx2sOeFY20LkUR8c7o+Km/3TvANdM6f854FizORdKUw1Csck9+pOQsZ
b/A5KFUPy1POeAGGNKDpjX9t5k8aRZV2VoTEy0qTLKSdE5gbKcw3RF/2AIP1Z1torSVxleqCeZuM
WT4kJmUvZOE3yKzS5MnaTEz7teeYvaQJhTuPhnK8jqtfDyo8pVX+3y0SvwZCvnXJbDUlETVW26yP
rr2ornT4+tHFA9vEdKaXOzMF7gayHiFWYJ5bAJyPbPXLEMtDpoA94y+8Sl+rse7jkqgUMy+ufkMf
maI55MYe6ZYk0aHyno9wNzskeygi6cD7JpUIY0Sha8yT9xCWaXOuyGHELhT1mr2NqBXQzD03KW6H
0RijYwg+UPm3Pjz28S278e8osKYT/EWI2SSlmqm3buCdYMhQ9kErIJV1Cuu5KmwU0BAkIkLTaJpH
AsUedyxa0sOp0GBX4nsVUc6q12yJRz93Fkb4RQyMt4mpZnx4CrjrFPqdRuHjxSgMeGKoEuCTnyhc
dLbTr24e88sPaasY/wlj8D8rzqzegv6xqtamM7LH0yfJYHGzZCRyd5TMrsKeDulj5QwUjGzawKQJ
LBq6gDVG0Oas+sqMJE5SguqDyzVsHZT2Ub2UHanbjJ6REGCV0ph+Gw6jmFQGV0U9omN7wgBOm042
sXs98CZanE3kSXra7gmrsGOWHVgsp3uURwajN47+2BHTuKiTX3J+B59UceQxC5kIZb1ezwnutV95
SOWXduicBbX+ia2+UR7Nq2FUwS/jypZS5KJ3n2qEp/SQ69mF9yAtn6rfzLb30cng1xCFiqpm+58q
j/7xWipkAqPgmOYQiPQQ9nbOEYG0xgtm2EVbdJ7lqMD0f92qjgQrYArlQbHdggQkkbrT/mIHK9jT
cXRZWZojVadZJqw7VaVNQxkgIm6FIlxGIm1DR/NVeABXkI9b3hYDcx0EAhP1jq769OoOru0MBWO6
lQ3gdFutwC13D3k4FaibnWpy34vzfC0Uwp7A4MTfgf8lhmK/Z8+y2LUBzmi4A3y29AMYJuCvOBbJ
ur8niqZAOUnOuA3jRuV6UuD+CRJAoFfJW9PB25cvuSIzsAsg1zxM9iw/2zhAYaB3VOX+lTepOx4W
ZImT7wBjXhnprbfPAtTkXM6AhvTeBWOsoM//d3bEnJUZFx3Lp7RPJrlHn9r4gY5nd0D2gBR1erMP
qh/6EbvmNmJiIIAg7Gtwuhxg97uysHs0RCxXKIJUYsD7PeYhLNDdXW7B26NMmAO4b3aRLWz9/PrA
yRJH2bkA8LK+YOojAkXcAKox+BhwAX5ohO9cpGOyaHTHP+1Zh7JnIUu7bVgX6GrjyyDcaUdx0ID6
PEGTDqSRyuijI+Ncc/QvLhiLoSnYfaCoKAvZ4cuixFrLAbeJoWxVIi5FLZ5Yj4vwMcga8UWfK1gp
g1QRdeAjVnUhgjTuerSZ2k8ScYML6SPU03oP8oStIEcqVl0b7ODsvp9VlUXjIuJSAkus5X+xhyjQ
L5/irnVO75KdVQQiFRiDrRlWcZpN+XjgqoSKYXdGGlr/5nu+xEKwE7juhbFIhZHZJtBb3rhrEb+L
EK7C9wf/m85GA3keENDUPhDQdMInLgPBdxjnDp5f+cVOAruDPAAxrGvYIhxejaRSc+XrnEg8pyP4
/6gIl13bdK8g16bFWzGK39eXFUU1PaiosiGqdhww4MuQ+Cb76/qBZRvsaQ3coG3YuwQ4+fNP6Zeg
iMwqsSeRoi+ANfLOaYuJqSvCkvflCo98XA9wTY88vVA32COGo01smiYNbwx34WDKOwmSdQhk2L8b
mfShmrPgoKECWRAbzTorfRUgNy4AU/zdEK3n0iwvLt4ZY5KoBUG+vVIld6y0O5l9rus8/mgVCJgt
YPCgt40l/vx7kGcp5st1rOjzOkUQGJzNVLqMXBrJRYP+2o+Dkl55tSlYz5lhLU1xEufhbcgRFbXv
d67qHAl5q55IlY54SEurbn4AEToO9IqVfFJHViDPgTOKRAr6OyjQPtNBOpCXmSCVUq5jyLT6pkXz
R2xOnJg5DVxQaGMH6OOn8G5Esolxl1ADkYQ/b7OuQil7R48U6T2BNoer3narz4DOqtohl1XBWJdS
IG1wPlbg0qsGCid2PB3fg8gXdBbW6W1WlLw0X6oRsH0I8PoIZr16DGf9sG8m3HM/MDA81gQAVnC0
FNfRVbGvIur8T//9oW5hMoZW3Yw3PZjD4jptABxnVdpH0hkOVwtlrXQHBfddH6a6OMoB+doi58FM
RrsRaklBuVSEOb1EvSdCtM+5pyB5o7yVIkAnx9UP/PXD5XaJJ8yUzfNSas3v+b2DHHmnpPi/uRRZ
ZP43XSOSNG0mClUjSEPeK6HsUvNXnmI0QPMBXtQ9w1slGIdXYtbMFdX0DPGqMl9kUtV4Qo2DWtte
6nFeh/cjPdh3uoJeifR/xFLcOoeKv88w/5UKYdW3myBhWGEgF8LO31BMYyQ1gr3jCs7OM/7cj08I
MAGqv45+g9/RdibUJnSqIfX2LzIAM6Rk39A0HnPZ3pi88J4JREd/4YKQBMNn4WiValoN9shSCut2
5bsMc09xfSum2sso/j2PrH4G8qJTTMHPN+wcMLg6HS3FEDk2p+sz/SeDvYwQks22fyL4PrBv4Wc4
OiKycDBCeaoc0eptlW2RNJEWEJk66qmARwnBaRq219xyarxRu0MYssNJbeaHmMWTZ/z9DJdUOFgj
lXTDD18ujMQjp99c4f8sPDFD6OSAqrHsujJY2MCniwlwESoJpZnGWy0cEhp3k4g9kXjNXOCTZ0NU
bmeEwuJvFWD4+LQEJKHA0rq9c+F73NoSyLaF1VsQZlUYWMGfElOqmv3hKkU/Z9p7JhGM9GAgmiHd
cYPUDYPgx+UZpA5nc8S39GB/delWotkNiakGo+PFJ925Dfmn6yWUkkGsAohvEt4U16FxfTnDETpz
+qOhFvMiV4dydjd8UxstUXYds3dev0eaUqJwmZRW8a3pj4afmgl7ZCktePWuav1p+/f+RLQsBq6H
IHMLhaOO1/ApapyDjDRnMsjuYG5dTy48p0kBXPkeAQruSq+6aElOzzCRHBoqQSmbpcK+38bkmkh/
ESnCddspOQPj2FRXqfMRbCBanLfUI4LywEnfsRJnBRnQU34gDRRvIL1KD22igTVB56eEPwC2pIox
cYn/CZjbtfssajrUbetePH73EgIaLYvGs2FZFDF/qLzV+yky1y26Flzms4GqAeys1E8zo0iq1tYk
72FSdlETAEflpw2jnWW+rjHvyNQQOOFxMqzToG1bHDCD4E+girSjspYre6nkPCYxeJ1TuSuGv4nF
rbIaAGGgMc8zvgTwzC68fLoz8T4QMLm88FwXFznluPtVn6gf7tyt/zgXfZG91TVGIcbQhDyj2dmZ
4oTLKE1wGDgL9Lj7LVD2Dvxa00t90Tx0K8t4oyeY8uxDi87rzYiFY7vhATkX8x9p4cmtV9fWUsCK
eKkaw37+2EJYnGFN9C+SSEXXslsCW5SOpUzt/9b40cAqUOj8+as8S6XhJlp/QNbykam7VDwPbV+L
EATmu/WGwbNhg7LdWzvYHvC4tT0zBQR3LeRZb2E2oik5KFGMffV3b89V0F2g91wlbD+ofp4XHRwO
E5T/0fZ9zmrjebz2zmnQpvL9jHQXsf0ajDzv4lpIPEKTDKJvpwsyQL8qWStPrkPARc1p/Xu7GBzz
F49QI68wrkgDINUN47K+KFNTLVrq+bAfZhpWOKJVDDmGMfRSBBN79uhpeTwDsTZNzMGEd58/hBNC
m2JNEnKK1w7hd+ZABoyYxrKWQ1nv/YS32cGm0J3q7pyzzUeuprS/fTn5s1M7QSKfEYFYG+nZghbY
bcqcpUVfnTIy0HzELISXgQdehZakzLGNhqzRUA5JpIeSL4lLF0n98/e+xvdeWNi7RYksjcLd0WmR
WQO3k0C3IhRXw/o4mMmOPScLgw4Hwo0V9mbNe+1QJfNsRM6n2n0vIUlW+rrffX4osb2EQrrTJz71
JAtvNhZ4ljMczbThPzZATTR2cXCp2OTzoxw17iS+jpDLNBECukVMBUg6ubUgr3l5GfTbHaU67OP8
mlBGQnr+LOvnBc7oXfEBCZyghLVMTdR4Fc/O7S1jvXDEQdFM/9oiResINuZRUsqDxxsH+rVd5qZa
3On+UPI+yjZrUi6qzN8mo2EKiYGnk0+fR0AQ5z1ARPO9RoNRrwdoqZwGtbobYPS+iyLbPPpMFeZG
m8Je5jrQLYKdt2TY/BFHo6moxcFEK+wuapBnhO1qn40FyJnG0L+Mj5vFHEm7yP1V56H9ALsMgYit
PVTiZXAU7Bz9lOm9JD2cogyFuMsSNMGoUYpR5zb50sD7VzzP3tnBvznQ9gnswJDpikfspQUG+PgE
j9lqHe+2lyDp+i7pe/szHvomSdOlqQOb3Dnf3Tvby7Z8B7n2eJBhT2eYSQPXaQTE7bq4uk7AM6R7
yl7d3Vy3VX1stA0tnSJm1n2c5zsZXwOyBj/PEcxUvEc2Wba1PEZGzJBvfjAjatsmOVRBzl/oTnqk
p3PqpAic7zvEliGRcu8yfwCjiIlJU8iTPnyhOih6Ri8saLbWCHPw8lJ0F4bTdzWQI0cPYMa4jDND
p+mCvHgfj+wU2nNh0tefN2oIfwi0yRDUq6mAkaJ6lPHD7GSibsSZEYPkRdcxT6PXOnyQytT0Ejw+
a8ilU/3eD9xX0BFA+3AJccwCS3XOkc50BxHQ8/U8mifPPqij9TeWL34W+sKMuq2M9jQwk9wQvZ+K
D7IQedqwryq9M37EZ9tQXG838T0wpMBY1Y1NWqnCLJ5kIFGR5LgDMG6+SUsCjRtWbVqSjgv0J4iG
yyWlnsQK83L8BPNKcjclfye3qp8BJ6rY7sQ5tEBEdbx5l2xUFa+OMdzCn7g28jKIHs9GPvu3Vs5r
htixhF7q7MPvJEZS1FYOT2XnSPeM5/ODOSfetOtMu9OkhyiNCZdv903lK+RA5U1r0J6pP0QSXH0K
7VhoUjR0or1b5nS3KlA2OoClqLoy65YiLuf+hN0ncGH+IfpbyYEcceHiYuAfKrIzKQ2HHw6R3YLL
37XRau0bZs2dhEPeM9SbwAgNrO3qUQn463oI84EiN+MN6WTuFmSSztQCmtzbuZEwUOu81H2pbUCm
WDWPZgp5eJW2fZs6/9UdBarGoLPcdbcXZ5P+5Cvq4f7tjZTWE9MVnZiXP5pkIZA1rNYs5ODcjNrN
2FtcBQC2b2++T2STOFoXxd/Yi1EduxAhva8oHEGrYWi2GG7sZKANet86WHqXr8ryYTY5wRSLgs/m
72zdSdpSakyQFSFZIx3cKd/VGAiRJxUidEcZ8Ry75E0wT+ZR9RtF1gyNOSDbRLJPBAI1f02cAEz9
pUOOC264/SHh1Lg9jmqUqXszpWOvHYyoQXBGGO4t9xfJEYq2pSHQjrOcMIzvbaDWdZ63GyZMhqQN
9qZIMOFgtrgtF80CgD9XVVew24ZRJgz87mQ3tW9Oq2vtoftiXPyXNpL9rFsPs/BeFj7Dpvr1pDeO
AryKe4SDrECRuCD3MnUMAbh7ndFAlMLUn8veKhqzUsELBb1bCljOHtBTqnOOFpwYOMCkqsqXt7jf
p20lCd+s02sVF4HJmSp8cYVZoWnPDVv/1pv426xqyWZ9oBVth89IRO+7EyMuKUaK0nebTdD4EVsA
bs2JM/ckAje/RLvIbeQ413zAf7sVvyOWvFoeIdjiDZeurujJoytAeHtTDux6YOtHwynanMGhVo93
VfSofUHqkV34JNLp4ohhAMOHzxtyRF854qqLNidK1ehuJ3sfRmi/dtjWeQmWdCbUr1Wh9ryWNPfc
PdsVgczE2rIzAJnn+9uyW9UkXNLWpHywfS6k/meLgT5+w0tKELfGlI2KW8Xbiaapbe+qqB9/AHjC
FB7Y/1kxj03PRtP1HoYe+lmPtFmyuBqrIjd3tOAs27sJriMFvB96JxJs+g8Y6ggsVilVYPtFMQa4
e090jKCVZkqyA5hAVuRbgSu2I1ydaR3Q3Ace3xu4DqAKBOmfQtGYElwAufsBDg6UowAdGWAUVQYa
oJ1iHJ0GbEX7cdNnyk2gDODz4r5hONtHohfR06Q1mAWBeFe96jylEBranocTN6SFtiIujzsD4Khg
/ZgYIR5cRFudOkYulww/GsCdvOZLDnackIgSHc+AQ2+zLDLBAzPoOXshFv9yYGz7ShJDmuOsbQo8
ZuLujvtghArOOHTOLXqzheDt67lBRP5JBreQ/y9cNjz9sOoYVRbo7YPng/ZQ7O2EC5uimD8iZoVi
/9dElXEak9B1T+4aIUltiZd/IywRYUEcs1pzhCoGishMCf0vl0f0Vxue6PgixhzSUB+37/km/UhR
657xcOGh04cNxWDP+s8vOfjd4izI6sYgnAcqTWZ9ImIR2fh5rnkfu4gLKbWejNaGiLmqccnTlDXo
c60VupIQRe8v97tOyEDZXO47w0rdSOKYXQ68Tdj62g3FJMggMcTu76WDlKSfV24nzbTInp7nnLFy
BDkp3S8WSNcqLkY20IwcerJIB9K8TdlsiDSGcRLE/XtDhVRrHsaqS4dwn0XZ+yLE675I4rhRYf30
2QBSLCaUkBoYS4wnxh/AkwimhiqQP6zzg/ohclA8afavkmfN5iFbkkRgsTJ/xzpHpjbQAT++No4+
heWfrI8WUfxpjZOc45uTylytFhS8+GKIGIiUcbGoKjo3xZPy9sd8Wm8g0LnyIr1tIqGj6IXmlB6o
TgGOkSBFyr7SyeE3RD8C4J2CeJyGu8jLlVY2kOa5V6KdeY1DnVzYzQbRlzEssqocDWwrxkNsP5vD
2ffbdpEoRr1s8oFihgILL3JPOmVYiGgB5eHDweGPS5EVyKY+v9VsmCbyXhFB1qzyYLqFMF+bY7vj
tP1+RWKEEkK4WhfJPwZAs3xlrAhUZ86Fgih2pQ5keTlSz/1qSd7xxmdL1UsiSr135rh66y6lbYA1
F1h8+q2X87Bee++wODWXerKZFKYkPobJBmYlPMEShLEwH0QmntgQFjEYEJVrfvX9/eyzOw3rj2ej
iVu/Kc8/2YWihK0JYdWLYbqGkEKQ7tbv1OWdDnUL3J2e/41KN65r7IlEH8bme8e81EYpEMndffHC
NKjrJUsGib2O409xrBKUY51VWffxgkRHdQqPunIlPHD7OPBKMxpE2MroknpbNepUnIvMgTS7x7M9
bMHR1AbxdUfrB8g/JMYlgl3S6PWQou22o+QPbPwH5eHJwD16jCvbs9v9nt4T4Jww5p6EMOScGive
Y7iOfSdOAhLoqtakFb7NmwA91IeQ2d/LUL1RzSkDIPG8b3ey935ndkHTjV+myLYIVjKcAzzphWfI
qiFPQrOWOog/6yaru1Rgl5TW42mSt2CgQ02lkltz7Nb4cRu7oZC7Y0tE6SXqEZOUGiJg0zbGpQn3
LdiE+svFKhzIvCqf33s/r61UQ3Rdx6/EmP7mcsJdGW4HxXGUgmkBlsgS9k/1NMvsh9C4bwkdSA1v
jh5kwrH53ncHL5596kT+iLo9jSpZCS9VbqplczPXuZ5sDLJd1Q2K5XfZCYoo5ytLM76rqqY7gPCz
TpMYK0V62i/53J0kRw070rcYk/gCXJl1pDyLuS+9FFkvv8ZB7drjRRhtB9tuly2e4Vt+yEix57GB
ZhOGzAgdO1DKYOnid7t2Guzxg582Vm3rpAOt+3qvygJr6gIggD7rtj56eOAcwQeVJeOzaoo54m8h
SE1MZAL/Wi4Bhpp+wnRP+Dfj9dTjPgcAj4DwxLVPs6wd6/NP6T+ExiIA7eYAmQLzjt+tAuNHHXQv
wRc2qeDfBeeVfbq0p9HUTcQgkPuRm1HdvR38kHV+L2O+hrGn6DSH2XcADAPR4kPUhoQZHJj5snZj
3JmANEdmjFwyYWtUL5fej6hjcn/2dNRDOz14IT4JqJWKb2Jv+DojN6jOYFv94R8ZxV7H4VgseOaa
+mIU+IJ9w80ZJ14d/F5apZoSo3gsopqZb7D0QTY/0NBoLZvJX+g3mwJXwThylWWhtDEzgU6GG7Q6
NKhtodcSw43aICgZB37RhrTUD1U2p4fPYdOEUUFPFnaIH5PaMsLiwduoj41WvjBLUWSPJDXe9+Bn
ffx6qGJRwrMEQQyF5QXuvbWY9bRX4N0MbaFqHHAD+AGkMCGk7erBlRCXM+GWQN8RQ1Cngxcro0mE
VVYZL+vEKy6tRmEdS2fn4UFdKmOrSD/6Dodcs8k25NDhv4Kg8IFLKI64q6C5kht3uZ8SdK8u/FLu
E7OppTfjdSZa60P14eWUFWggOcYbG2AUV9A/Jsx6AMLawjxgY+yKqpUrk2O+uCriTJnCgt2iIYd5
FTU98OG8mvmb0iASeeLDLYcQiVM7vGbwr4CEZexCdAPgqESw6ez8izaBIoWuNXT+RlR3HfQVJu5/
/9Se6gDDTw9gWzvhKFbmKPGQCcvT4Oqg/tXUpjDzOvir9nSMkItx9fVXV+yeq4IbQ6+aUIzoHnaQ
oZk1hX32TbZ1G/iZ8gPomVBKX6IQ+3eWH6HyPrNtSm/KBLkZK1AMbSTgA4mjrAIVYVLbRgUPQ/QR
leo7hdJpMdjzs/LayeSiEvUCQR1HeQUkA07XxLRcrUkeJhUhfghJbhgbLBd+Ovo4PZQ8I2theN7a
gS/U9llNIQS3Eer4i1rcFPLPuBkvQCdVAxuXn3XPvgO6N0ZXFbhi3DBZWGh3kttIASoOsE5MEegm
jJpDDufUDaWPFiZBxh6y0RSoVmSm/PbmMLh/2sWBodde6jS62LEPA+iewvZPGrYxCTT+19iCrXXz
DLxWs5wkRlouWPzT90zZS1s+dYOIsbuMLrQVxnTDonzDLKuy3kbB4TacUOq9RxjdbqudG3NLL//P
z/aLzvKyNNC4ew8ZuQG7n8kUoymyWcSZB8vVZmWm8EfvzygHHeUxK5QVyq0f9qR4Gb8Qt/PXDL6e
z37HkN4kfn+Lxfobl3PYrvoQqj8ycksdKAijw5TkmGgFSi5dDU8zVuQZTVXN1e6dGDpIpb+hvz1e
+WsTn7Wjy6aDZoHP2mjdNEqDQzj0L+uRdWXHBW6dRJOE4g9G47o5YWJAZMpMVjxPVITyzqNXUDvH
dWQlVEciB/SDNX5/+atzpsKWGMk4xTU9w/oVRei8bWOh/K8s3X6/xBvjJfoU0FDgGVdj3FTCBoC3
6kLsR7nsjigeujoJsGAKrPeJYSESzznxbHD2F0lmw4stQ1PBcWxHCfCBJzLSjS2V3XEqe0CNDULk
ZxWYgUBm8OivSfn1gW4J9ju+VrjJHVzaIPW7EGrElRsoxl3EIUOVfzZEEZJiw7LgPgKeWy2jj5NX
DpUeXsGb0q8l1hAOm/zBWFNx1YvCI8GwaduXpTpKvaf9eNjCgc7+1Ia/Mcs9EXgbIgKZKxrrj//Y
ZkL1MKgVzf1uF1uc3a3w1HmYUa6NScHI0Fck54M+LGi7cZVJ7FKcYx+tsEB2QADOw3H09pg52hiy
aOgpJyJIc7HTvjidmKHflmEZr/fvTp4Y2xhlWg4hdWyjsSzwuk2DxPUTm7lNxnnIHbU87lqmOcUu
YI0LKqYhtwceTn4NVZH8dZnzrCyvpKezfRxUVsmi/FxvZsB+NqJ6t64Ib2JcAXJIf1G1RpdiPG9f
dxKzn0Ew2u5XK0csqPdFxG6l/T4EclDC7dm+eROdikwImZnWBoPmyI1/Ct1cq+JR7BAcn3ClsJ1c
X/ucGcey7nKJen9J502w4G/SRth5f6eDxIKSbcCTH36wompVNCwINdPdsnOVXBw5nS6RZVu53V0S
25DyvEdBptZbia9Kcrm67lYKWGLFVwcwbi7c+GIvO7LbRXG2bDP937A5FWdL0hrDoAWS55EfhzFc
mhoS88PwdOrQRZPaWOpg9Ezw7ULl+IRRnpypqCbr+MpRwfuCSKCq9xhbGwTPihB63OgZOGo78Fqc
7+BM0U6jhaYvm9ZkOJ/0Vijpovo4xuCm7mQGHdFo5RMgLeJ7Xc1fwvsVUjPCWMqUEc5eoIzzL3pb
2YanqOEmYnuhqdgCpNJjF+FVvd7qW+lXeQTupP/UfnWr0zrnqUMY8ywizFTy+zurJdfzweHHAnA2
eIWb0m28yZ/7O+W0Ihho5yrtKttpyXanMU9OJ1GOhQZz2B7qoMci59kjLtAuUYuAf+0rvzG8dRq8
Fs7RHm7YV5OPC8kSJI8IF5c1ZO540RAZXMJsPID1nTjqmG0hpFsMXQcdUoq/AmvncWALpojJL4xT
hWFjmw0wHvFALxfrB4VLN6BuJPqGJO9WPXlAvPH72Fxo/f4/swf8O+I605UGiHbNV35+5+I+lRNf
9rdyVcQWyT9flDuBE5IrOCHdsfib9MHCals/Io+aOCbR1l75iH6YurdlqbkuHhM52VTbpSA7WdLB
TH4NntMBvGhirifAzeVtQVwpHfQJMq/yAUiKf1IIPWIkqqf7Hdr1b11azq/RiyWDmWb39NlOx6Xh
H8E1a78AxXRZm1x++TchSDNCpJKIDK+HdVwwhUD+f6vkXEWWoMgqt45SEwIhMf8l6vOBVwkVyc/r
zcJ6kgVcWGbfXAl7N8uHRQtCEPoPKoPj+kojXbnthCHT8RWWmVYu9ARD+gZfw4VofxvzCmSwfLEr
ePBWh9I5tQdK59IH0rNMpeKPZfi5ag9EjTBmQKreHk4Q6qOrSlBf5eFNIELuNVqUvBk/1D+ny5aE
N/QAzor4DnCl2oK/JL/mEi23pxBTPEd4rHl1tFjg5Wn87DTroNENRzEKJ+6yU8eaKZFDnnZOktoY
HUeGCM2p1iH1oWE61RLxTY/FDizgfc3rWakbd1uieLEBM7+BKQFLR4wqC+TO8kute5hvB1GxQiHx
3hemFfhtBdcRVQ7CNHT19YyT7pPui9Nsnk3HGBUKNaGbzH/fed1WYDGrqInGkxE84rioNxPaM+MQ
OY7DF1egarUEJG0NvpO4fL2C2LweLg6oDdXbyZEfE5dxh/HKOueYHUGeR5S913828B3vbHH2ummN
VroaoHs1mOJCp1BKLwZiCsMBeGy8xbX65a4RWZfthevxa7AJvQxY6sDUOIhr/ZK4Mlp69tojwVZt
a47k8RY+MjB5gFPYrxH1pW91hIZHG/0Xl7mrMXXbocLhbCLZRBPvEyLA3KHG/3/2fzyOlYXn1t0Y
GzGHi2ptBe1MszaI7mpA6WYfu98Wrv4a818AtnDmBUt3NbaWmHP9N0M/QVNtsdTz5PqXShPJAeS4
vgRVQmx25bNLZBhd/4GMwOcsdOvFzBdrL/WBccXFTFhqFQBj9q8suXXXwedDGvKe5E+mlTLmCEdC
MXQyHKWIqcTuEmeW9/TBoX1RBoTA/f/ifx+9vwzlrzKPMG824n3bGGt/RYJ9tbbV3/my2mTi4foG
67POp0Bf4wFpjZJlQEKo17rXpMlJsuK5MID8ViADup3XI1cIlW6Ex1Rnqcz5BFKXvkmzU/6ON2Na
CHtse0Y96oMYXsKPD0r5fL9ctakwqxDkGJyHpVsRvejk5F4gzEzY+r006xj6aKT5unpLmjqEapsq
5ZuHHDC7Ddzu8kRzpnIJjFxPXs5O+ZjPxiVycEf4a769vtKkVQrpAPJtGkYRa6yawmv/Jc0k+uH6
SDVpj+AJ8WVKJ4QPHpq05PV7u5LFRuVP4Prtap1EsIO3iIH6PP7MeRC0ER+sa3UUNMOy1ZDCxDmx
D1yn8mAjbW/8nvXoanhNyPdwMEUHJu/75R5P64SCJm0dTNZZTmqzeW3XbFiJjljhJmIKaa5GojE3
x/yFBY4EQTdN1Pw62jjhKbo6WivAaTcrpx+OFmsCTb7hnR0bUDxn5EW51iPdLRhEJr2UgCaudDk+
/o4E8VyS2f9UAkfliScWCJou6/bQryyJFZbj9dK9oul17sfkY7UktzBfNNQyRUuFaP0T/kxanUY4
DVjeykvf7LU2iwEfnLKjWbgcr4KzjsRdi0bFkUaFj9dZ8DEO5cpnX/bT+eEGie0oc/FMNbQPwURc
GioXJOJpP3jDnMrxInj94oA4D6n7+eUjMIgLU4QjmnUMsFU2LrPHkGeDwD56w6dey9rPQbteeRir
3TPaAEiOiLUvblS9SEBdwB0Tqnt/kXQEiOcJIOTT7t8B7gaINHA2MoBbveoOoycnGjmlDVeSS/7E
u3bP7x4/PupxOQ54hr/RyVNTE/qsRq0ATIJCstOeP94CAqaIxwCjlbetQ1OwYDTLJJEbmYwCrp++
dCLosl+99BIUuButuHEF0hSAZCQ0Yj4tBN691c2wfnji3mxh7dqUBaya02AfahDsh3KidWJ5qh6f
ju+7lKJ9Dq/qiYIWfo826qOAngXBF34kQXhmrKF5QFpSVzHpw/a5x+qea8fRDrufzdomIbakxJhQ
v9gkg/7/bI6EO68mEHOkm4oT84Sass4reHTwfXyAxDEpkuMVAz0JyNZfLvFuIperk2Mt/bEfmOJS
cWHxIXMUNOfwW93OMzidUxhiJYSsdyB0omS2F8EnG1hWx76BHETinpeyl4GPU8z/HOlpSsvBDKaV
h3rhNh0PIFHTsbgXtJHYnOZGhSEdKFXLEe73lGQ2aT3/Oj23yW6iele1GS6QbanocxNDdHCy+ZhZ
wUbKvpk4IHqZyL6cOzrKLc6/2SMLLccd4wixixmE4GkI1clncgeJ6qixjVJbXr9xEiBnVVpwwWjU
dlFhV2VfsTorrmFNi1dfH5CEIUe+wBqOi7H6Kn/zsRIU1hWDbX9ZMSH/I5bvpg03MPoKust9fhvn
KtjmWtYyGa7FU+Lsandd/1q1hZN6B+nt54CrZzYEBgdjW/coXMijGFimjFvPYGKqbHBXxEkjXKjL
ktl7U/d9C+L9CARmWntW4Ffjq93VU0rwnntkbEolvBm59L5q/Yw4LndXKBqhX6UQeKHQUBDqepnr
v0Msfkzv9F3JYj3fhUMWvUaTag9pFDbh09jO08XKobU/asb9UYQM91sRKO1wwm97RJW+7bspG5lJ
CvtkYcOBvdurwA3oVkIX42LDxlc3AabqNIJbxDUuYdyFWj0D1T71oCzGJbNqGlWcQbIMAr7onbdm
qB7BhahEo80siDlKaf/+LDHpDoVGYds8vW2qlSNMQ3SZJXmvn1/N7L2/NttOn35ZV/Dx4BXKRSF6
RxdjHHcHE6LSRhCAyYS9WtQUwIwQBKBZG4pvUD9LDMXOp8LX8MVlifmIlOZYvYhTQoTeQmO5vg6K
Uu4chDu+6x5DKIsX/uSJsPlqswIf9g8HcbvQa45c4pNXwcLkyLFfTyeWmbP0HAeCWMS0furC7UFG
JR3qHMNRQpUu9Sd5ieMJdp2FKx2MRtGVxP0lDN1MC5iOOJrUwxQW9WPYkVif0RST/pFYrfo98Oa7
r7MR+5ZsqyocFaOwRGAPLiSfWMVx3PwgNUw8PQ00dzNqGlLZS80Xwc2DCleTIr7W1bvZY2bFLcmX
xVMFbHY09FpsmfAMJoXYqq/V3cEZh/WLG5rXLBbKZVdFWvnOzFLZElaEZ/4PNBsH1h8tXjK1OT38
1Fo92hYUEV8w7oUIBh5BwL3MsyZN9y6Y3JX8MKysO7vXfgBMZMwPkIDvs4V2Le4WeVmUNlEFrNHX
tfCKajmqjPdUHi4BxyJ25Nopezg7fUIm4WV1Co+I1c3rLzYlaXos6umRE0UBuCdYbfxScYuynypC
piRhwyK3b6uW18VvIo3wUJDjwZVc1CFu3TeH0n1OpkfJKvh4IrxeWcXRyxUsO7GTgsI2dF8WfE8Q
PV0uxLzigfWxxdmRBpYJrI/lRjmBv2IOjzgcwdp4RF6H0RMlnlmF9U1L59yYSV1uBw4sKhSmbJ/V
HaHi0GoBkEj9H/Iiy/JORqp+w4XSNNdj2kVzmkh9p//7Nx5ktuERfoTI5JpnGp9M8umU1dLvzxRu
A4ABUT2BuAXOUqXU7hjKN11a1ImrfwaKL1fNx5bC+0hU7MtHPCzk1fED8aZY5oTa4rIvPpzozNNE
+gzC41FEVs9GGeNzxhGGGLMSxDknqaN9qOsltHLfR/+no10iKPSA06mq/2qfdQ7h3eR0wbJR4dg8
FUhpuygZFk0V5uurmjgM7oKRbT8VCm075tS44jW7TCqlTRCXM7IpVWJ5ceOyDqa2cCVOSdp26P7Y
Xe2nUm2WoldAKGYpXBD+GaTQDiS5dmGnd+oLxuzjEpETEDgInorIJgQ3Mh7IPtR8slET38kH+8tp
McLu+2k4eraXzBkrCNw8ENQrJjxsioXV3eXEUwcjdIn7DBxZ/ZIlC99N2w2rqWXtAcpuqkHGV8Ur
Eh4BWTA3fMdQKwhko/jRH0/yyiCF7XgBXsEK6RrQCgMxkfD0J+/7ZZTtZkOeuvrI7QcjMSIeddpd
SEFiqjPzaxTk96rm/JqT+YrAHEX0LlFZ78/yZM8kRs0Q1yoW+rQlPfio5fErro/Bi0vISoznkR9/
l93mzkPHlyj/iZLVEAD8Mydk7uEEQ4ltSDExIt4ja3O756XGSzsg3NIIhKxaiq3uwD3944USY8xn
BrDgKvXSFDZKXqJwpUjtVdpOxfyBeGG9xkb2SJtpDxDx+BjRL7DGjMpbnA8Vr9UlZZzTs4LnOYx7
+MuB8Zx9vl3F+jW/K9my82EvIENroEcPp99r4rkBlnqf+GtdQOvw24O4KjgjPAynXtOu3ZRVyXuQ
Lfbb1oyZjW3GJ8R4OIdNvrlkhv1U/Pn5OKiwRrv3VM/zjjfGwyAFraXX7+h57/9oeCAzakIRwA1/
FIoWQOExYSOv7q8USqHVwrB4yVtL7Zrj3TplzmJPk4X5IlJ9jZXHrpE6TX6Vk/iVkC+7LQvggBnr
IW/CyUP3H+kkqJiAq70NP8+PvDbmePwVy2+R2788NPOXaiuSzMxB5LdMMETQ74iEqUOvMDZ45mME
z9i5xMMLRvN3a1O46O+Q0Drod/BZ9ZPj7HplEcPY4slRTZ798eUe64rw8HsVl7scClvO0pDKtJit
3V6iJw6UiRxT5KV3UAO+Z31dI9as9QH0Z3cPchoDmk+X8dgwgzeUWcsva+2MTnIlDOR/sxmgaDdP
JYYjiooF3h0Wxro4QY1hg7YS94xQG6a0oehI0zU/eS/iLJMIeWARG7OhUXOAHL7ba+CUvEroKEpt
O9PuDUW0GZz8OViDLLZ/JO0qFqQwh2VFo5ulRtlDpbvEeKm8VBEXSc3PEQN/9g0N64L6Z9HbBO+/
j/b/qv/+8//QeWPSGuFjfNmO9hmPs904KPyMZCTWZSaC1k15Nk8nuz9rMbCx+f9SCiYr/Tu7SDS7
EBbW3Pb0Ic9uwPVlxGovnU25aCfrwO/sAoaDLOXyAUczob2roJOem0bI2/WoyfJJNcL34WOxP0Tv
zZ2QBDW5nOvEK8nUMgpdPzFJFIWqAlDbhmWHUDVcqKihjWerRz9YuO/vKgcjfgXUQECzGQJuOLUs
DJGJXNkGx1PYEoLkweau2HMcuEw4xc/rBEJg2k/qmD9R3BcWJRSFm8hWTjkyPsvPJqGxmK7YBsek
YkUB8FPPUWadL325CzwSq7EZtQHZ4dyCovx+ST+ywvp2jJdc+6oRZTdWRpPHmdMhxgIniMurHyls
/uoR5OlzZQt8ZsRh2tjNRh4f6PmfEDJDsriqmJilBp/MYQo3vHpCN1rgQ1sOKRNQ/QfKr/zdDWaG
Kah7DdckPgM6cP0PrChJK2sqxoTFeHzg5tRwIZ0xkcGkPBIa/TNdJpMADjvcvcxu8XR1UQbDJbf3
JDy5XWcvJ0/J0YtMbGqMcHD70lR62X00/4HLbjK9hlze207luJzEDahYI91c9je8lNfFPqJMwW+K
pZBHj5y1NkWkGinh1TGw1uQOKwRBzGKZojcTOSspl3f8+tP+YcaL+6OnmoZ5fz/BIVdTBP0xdoUS
N8muGamtKIVeAAUrIaySOhGvUIBR6cZeo8yO2SNjyVLLyRMw9OgRZ6MVlfg/Hga+AnaQkWm0YdQu
0SwLHlfcoq4inGMZDYkRashMHGa6XBcgLUc8p7xvHlC9jqaHxA1fUxacBUw+t16WB054Yue9VRyw
EWjGshhJsWZ3qFW2+eZZZ+BDG/xPXzPvPMa4NX9C74mLFsVbDB3hR5JPJp+210XiuTzi3IFWjyNP
HWNVtpf1kUr42WYn8s01w9nWKby9K23MB8v3MeqOsvMRlqr3377dlYx8DTCNJVCscd/v+6rzNGUW
VW1Hr3ZzCL3EgSsifqvmGmp6FQmz8TJDjFvZKrNN7sW8WHCjCsxgrxuoMjpWYIdduCyEjolymaAF
m+tx9rkGvuwOvlu+nKIHj3g5WyXDYlVm3Z1jXq/NqlJQkxX08ee6iGqq1K99iMhNcEH8K3yCi36G
j6kSx73aH9nwXPMJBtLDqCPz3ls/6lbxIlho4HV7E+0PWJCnR0VJe/G7UwaOMGP1U0+M+h35b02m
IMnr1Q+3uIRwqiErMAf69W5ktPVazg6v24DQHHPK2z7NGkxOZQ/EbEnuE45QsbK5kVZi+SsGUxg6
BFaT3NPx4wefB550LFdAiXLWozz6JNhIcyjnG9+mQU4InGTAPbFEecuL2hOlAkU0qvNDm8EOMt05
uPX0IDRHGWVWcq79y0HWgEAxYqW3udTha4XptAvmodeCun3xi9zDHdzfidSdFpVshVIAu//HyK7F
qBktGTF1SGcB7Iu6cjn5Yl92JirdNqNm2Xs8+9Ppe2PAPYRANbfIkHfVRYWN4bYHXd/w4Pu4xGO8
GDh/88nRMgUFKhlRPv7eX/kVU0Xy9HXfbHhHoxj2UPCkPahsAZAFSt4u5FVYsDCmCbce/nTmIaYs
bdctHrUtPcsEzPOMgy5zhATQDnuSH53+ZdF+QZYzcte6MVzkFj4ROKI9UUlkdeEC79EI4soqrsaJ
86ADropqDEzXfI1l8BEW9z907fdUQNjgq9R6NHnmn/BDRqYll8ZoTy1JKewErd8W/qgngnO+gQrm
0WX0E0J77tyuytML3E0QGF7W9Eoh8V5e9Hj9G45rwih9s3eXmzTfBQb/4MF1puhLQbrURmeew/Xn
37vrgKlcJLOEJYigOVjDcAGs4eEHZKcVPYpngcGglH3y5uSB/nsvf2WA85OcHJY7MSIum9ue3T6F
4h8VNNDc1QaMFmur/OMBblJLznku0mM4hMlsXblnFCpGv+xjMMoco75Zs838NFLEzkfHWV/c3RSg
ZVhZ7T0wPpyHK3N5Qr/DR6sP8CGyvTmI/kr98iM/jMpThQzhEnk3xW+x6ishAB71vCYe/OibZUEK
DF0+Lhil6jrONWErYLu/d2dD6VJKa2GkXg6+Wqwl86MKsGdobvBXSskfCBhpCE7oJcHpmutTWfbv
QwEKn6MHvp2WXpxC/blIa0dKxAlGDu2CoXoOX5s9J6mQac+zFikKUGQImqBPVPYL8gXl6zTMXkSs
8GNM3EaNaS2ArTVpSqdwDYS5F0NYizZBjF0cgW/93kVkZvttuWiZ+oxetiatOIArOtV+ovQ7wYZS
RqoPNnQEgvRwfvIGmC9zE4MWF/mhwapHre5Nuzzslpw5K+8BlWyHYNc2a745/IVuEoAVQuGaBLeT
7OVp8I9uq5Vtjmx4AOFONOgJJe1Wdv34mhn3BfeKDQKI8yHV2B8mcRUDwUJpMs3S4anfcKvDr9sY
DIaiYSM5HVhc699RfvVcw2vedAkZzIZ6DIvMO50KlCfyr+3p6Z6HnzBG/s9w2SUYZF3bZG/K2Q3W
nrQpo7Y4MV7gbexm++ZojrnRn5RCks/VNg6aGF1q3MW3WnUCin9bLIeyep/bZUF0ATzsGSOf6AsX
JjYXeEtyP41T/13zzZsv6q8D+Wr8hUwWzQTfrL/Dpo1GWMXgFrx0/YHOs3g9bjU1WLu2AD84PA/q
VE0pahsgJsGZRLtZplZdRXCaHO0xoUpvCANDQMPbKYYZ9p4py3+J8679HyKinfZOaQdbdSVcH3M7
Jc594hfhJe59KNwSRyUIsBUkoqsXeCsEIkxLSsJ4ca15VwU39FnSHoNRw3l2eKIBQAfZ1rJvrbfU
1xzkVW/6Vtv0pfA0sRAlPetYlC1bSzNzfIE9a1kRCWYr7KxrDUs2GKpxvO69fcUugvOnzK471yvf
J9UHIQiVWW7tw59Hp5tVKp+auPUE6PeKjacI8/rajVkstRhwqAVE2q3J4RLatCDuxHXUE9+pWs27
mnlpT6/jQdrj19W++XUCDsk/cIpQ0DaLAKwyCD7EA8MhMzMz+vsN/yaN09kNZ5siAZ0mKpEw4zC+
2GGhesqx4poXbKPfdrbrWXn4HM1MMlM8p2Lm3NPly7+M43LkivqxpyVvZyIym2uRABBZ0cna4t2T
UDLDZJl6SPxS3twSgnKIghdf8TirJKJc0+ALY9fR3zG7ffihYOjH+kPjuXP0550p4S/y5an7pq37
HuEHTm+kRq2Grr2O6xaKfzFQbBUQxPH005LGSHQcUvUHUlezyDb5CQWgWtUCYLeCLBDlNRiESDLH
1NIb7qPfHHtbcMFd/tmE90B3s+2mbtwPvwABry720G9HpJ2F0/m6Am55DPlU99tcbvcR1LBbXQma
CPTdqlQw4e9MhQuHO9M9j0bc/htphHSBHqmIkYq54Pq0VROZ+fV5ocYVZ81W+NLLalbi5a3VoLZd
DmWh1mT7dSs+tVkJm32Pql2obnXKNXaiXvfPISKU4x8yutPlgKlXr3fNdu1zcpmorwLYbSLuf9Ky
vibdrdilDyZRzYKhgPTmtBNRIcSJG8mKQIsizYghU4XS/pKbxryu8PbvXqutsWUx3njE8EZiQDPJ
izn+lD0ZlOXyW0Dy0b9E96UQZeCpJMcEKHcKcEyHC3QwWUana4msY6AExkSUPWM+u3myLwk2Hvmh
7EbS+6s707ERg5jipfW4Ws4x980vs2SKWEBqRyhiVUZ+E50mN/Wm9WbVSl7s6kw54j9K5tuIzQp7
f+CFnhh0WlA5aKotNlFpGfevg8fTWYqFrT/W3mH6roZR1juplq8/GBVYZYobRQqcp8GmO4TRixTM
qlWp2/xjoEd8rFGWZSQZ5GtHbwXUquM4yeTkcdW6P0n0AdQhOAVD+vBRWG+gbVeh/IEv9gWsqyUw
GnsyCL58wLNfp/vT+mmuqfYKI/MVLzl5rkpxbSyhtd2XbKzKo1n97+ymtgo8hUzqZbSCQ7frEjLe
Z4XpuPiBuGAfCuiRXHCxtcYd8gyMm3GGM5mopUQK6XrBnWLekBvjxyQG0fgtfAdbRMyCcYiL1x1g
Qbp+UHkvSIACNSIODR0mT/76Q3ItUznF/QS62jBCMvWtovNBTM6lwLc4Tw5pMenIykbTC44aso2w
UaOhXaOmDDnHHVP/Yt//i0w0BGlzDIc5HwvjJObaRP7k8EI2lnxfuyez8+JvEebnxb8SVVwbubGg
1KR+zLIdKBCK9/AUfR5rLVxFx1KAhLE/YOpUoX03N1nrb4ddeMSQEjUaEzuuooLrruvdB0KrflgQ
KFBbEFMS/t0NnYEP4eSUVhYRuFPXyczSv8x45cgPqaqH82E7cAdBGOcMieiJAoUmKgzTmi91kQIi
9XQLqxoBv6sJTXsdu0bhsNWKAxX8CJ44lxxEqtG974b1CQaQISQS4Wslxtl7ZgA9vCoTShZdqr3i
ZvQyreT2GJqAo5I+unH5iRv53p3/02wyQLIzgYixxINk6fyPUa+NtRCY1UWgR6Sh8Ws9tYjgbpL3
XMUy3gs0GpT5vlcJ+y310ZaoRMPoNmFOTAf/SAFnnwH/HRrW35BGGLqEm8GXLCTlrA3DV7/kmoYB
rCqzgZ6OocvhzKN0x/iOFjSunlteN0nSyUHX0cu89lAFn1hi47jpH+bbgbGsyFBiMRDOMuDCUfLG
WWCJByyx0QG9MpBmo64rtzd2LT+oPvP6fAAH20BvQHfPormnT2t6puch5saZqNZUb15HMUGZ5OUv
ce8zIQWoXX8jKFlP2Nl9qZ3r5QZSJ0SmqvdqjhsYerbypl/5RZTRVUd0RASWWnQ42d0bYbx5kPCW
bj04lF3+nJZXcsOfilXjAsmtSHMEuxbZ7/yem6WLUUi0KwKPciva9Vn1qb0FDUKKshGkC/AYH7O6
m93OWY4dt6Yla/LFTiSBSfjVQsEKCIVTTebYnR2rnuqy8HnzaD9/c+ocLFc2dT7h72d5a8wweP1q
RLDusYHpfYw0ys4LJJTJs/dmfgd1E5Mj24HDPK0JYIEaBctUMoBH4XqpJAnVoVUoCptxMjKLdCb4
/XLbOUtoiOeW7d94uMgtPoobzr36dmr4KEQwCXKYsHTochKRZzVCcKEOi0zL7m7EKZNJ70Ju5wCg
W5WKx1MHpUUN3YwLfHS2SIDvJscnNjAkDd/tm/6YeoTBK2sCqw98BtImFh2YeSCHMpVOr5B3lww7
29wchOsZbeVB1CzTZG6i++OAtFs379UAx+EfX4fqfrSwvSsyRuiqxHqcBSRwej3Y9h9zQjh5G6L/
+mkYEMwSvHSQCffHdmukn3opPlVDbtffZCg3J01D78ZN+GTPAJntPpF7RiyW1Rhj+RiyDjXYs+7u
Ne9ISzfibZcI8Zq9Hj9b19tDkvHmd1+8PrSBOlA5jrV6Pw0T7DOb4c+LiRkWHUXyydGTYyS95Wjy
x4ul+kOK5Y3swZTJV8T0zMAQTII9PjkvYfQC1pMO6wVzljTcLWAUohHZi57kEkF3fHeQtgazPGdB
eeBDJ6lGu394wM0y93jOXBd9Z8VQ9qoMVXuBFXXOFlv8LNGlXON9pPpD+J+EBB4dY2tL4iBzGgVb
2DfnwVDQgJ3GnSYql3DvikfnyFGvO4SfPNYUg5WjJmGTxbAdVLHjlV4eeCavpKr1knG3BnCu7wFb
XYxenEYrpdM/DaCbMmtZFwD/DuGu7OQl2TNjOOHIGMQoe7uDjKiyAhjXsubJX91WkBCQJwiG+Ni4
gSp392hnP1Z4lr+HpO/DisYcCjEvzm/mmDr9rsPk03Nxcuzoi7druEnZdf39oyGwIauDw/qSLE1Q
Q3nhHSzhUGFm+v5ZfVkU1OMhZymZhNbF6tFjUoS6bjd8SvUk8kWxLaon+UHXOUV45uTVF6WaZXOn
qUrqTHR7N6kKbjwUMZNbK4Q0psA5b4Vr8okF4j2myDEl1ssDgusf43GYBhxlOVNs7DI9vURhfXYP
7leEwGZoDgi50wEyt4Up0Ep6GgNB53BOkwkQKFuiYu1B7R+MMikE+0ioozxkzn8zETKoyMx77Yjk
yQ241KIXC5Y+h4V4Q4+SRN7YEW+FHR2DWdytkoXOcFypHyfsswiPjR6QkOQGK7R19/CV7U/p4/Ql
egAscHJn3hsgNU2/X6GhotrskaS9GaDgSxn9r2l+W1Y7oUDSZlmjDg3Smi1o4CLS+6vc+QvltdIJ
2jYmEvMXHi5S4q5HYNuWYHgfJcqbGkRF0bQSMVucz22gvmvNhFPQV/JFX93RJ+PJta+DXywk3MMm
/Jg+j74MJ4xIaoQHxCXa2FAynVRPRQzdmQ7e8+VIq1l4os/jO2IPNDHS1HYbNzntGmn3Oy24mTl3
urFCt8krzJ2VHHthAhybz3pVsj3rIfqZBJS4zmvmKNMChbkUc/FohAIq5lsRQ4mydV0zjTLZKW2M
zSGb0BfIgssp5HNa6Xll4gTv7G1AF76QkgAjYHWVab6a2Y9nGtaDX+2atwTtAwAgUomRw8cH/xwV
JyjVdrZO1AzpE91bchoHWM183AZ6SyNZEO+GvEy+Zevx7m5dQbO+dloxO6cW6BIcC8LBJTVvp9SB
UVHSoku9SPus6th6ukmKVdQsA9o3WP0ZWrGCNfNx0dd5QVMMIOpTI/UhYEKyl42kqay1DpC7+/v8
8OyhgoVqymn60lyvfp9zYXqtdxjslzL6Z0vDLmgU0trKWSYKWF6ct7i8uQGXDo+jh38USu+5ufQR
vAxyFpPTx79Yd7vYKn5PGvLfHU0zb1nj7WAJERTEo2eE1/beZDUyaqGoMcpXQ31w+EGu2T/fOpo3
S3WcVjG2GI48SgMceGqSpcxDiUpzDD9zBGk8IaEtx6tJGhaq4Wl3VGTpaHJOjOlQE8K6rDNZT280
9od/zqr6NgarjaQ8ehmS4aMnLRdqozfsX3/Bawef/8zOVE1AxtltqCG9CkPb3breCP+sBHSvVLps
iMkLfNJbaBqOB6UgyqCXwY09Q2bIXoDZrGLMMCmI2DKHLNDf9NwBFkFZyppnduAZnsF7+BD3QCbl
bTC55q2/6WUCN3xU8a7uRUIeIUbi7DSh4opBoCcSl38YV/fuoDi1sYfkNBl9w7XZLuGX8Zqi8Al4
XpS5i4dDE2qFurOz9bqduzp8xJpOWHGImwf1/6TfN1D0tlhtYyPcr36RTuz5khNv1Qe+TvhfNe7y
wJctcfsticv96cS6GlL0H50MGz+JEKfnEYmmLMdb/Ny1oYXl05GyDuDtLjA11rQ59t2a703oe61w
XEy/Yr5r6W3DrniGGuuLZLoBxX6W/tll6SBokAABIB+I30yPMHjiKq5z74bBtLgwKkrc7HMBR0vt
Hth1w/QVtKZOR51Ej9CuWWCbgBD5x5jTYemjuA37ugAWKthoZi2eLb7rzyqwVcpsY3P1p5TMIBtt
WtRdlSWaIuOiv9mn+ENMAxfQb/L4YKA/ZfUywS3b5ThVAEr2Zj6v/pnrrg6jBTWLpuNyiKEahCsN
L/bi7EEljsOmSMJEV9QVmIEFvzNd/2E/Aoei9oQJ0spGdajUEPWow4YN3DLR40OveqKwsXABWpns
KBi65igTXCO+aokrxabURuO0B0QcOg0W6CXp0gOoOmKw6B3cXa/1IC/vZ1RQ2vWqoCytBEGNWl7u
b53fpqALCTu7Wz38KBajUFkMmxECE8dQ5tAXlaJIpMjAzUiS2bQxCFBhwvSK/iEhkbysPm7BxUtn
1qHyZ4RNBpBZvTIGdl4xgiIkUxRGBg2W/7vtOxlVIUgk8MbU+pzw/3AfJ40UeFO2qxnjqshP6Bj2
X9Y+EPeLdDWUSe99c/blBjN5j+uU+Z0TrvwzceksbNTqcyId5pNS8/TqjDbBufaxTyxJE4pl5VMB
bYo5pm/wIItx/kD1Fe5aNJCTLE2q7gQCFli+MfgLd6cye26H1YG7YdmY+xw7yqy/6Tc5n8OaRkL2
96T4aWzMtU4eGCZRd5pRTF8uCRFL5watKtY0oRzWeylMqiwe3QltGA810hvhfgMIWeX3ofF+nY+m
6cs/MmZEpwvC2qUmVK+fksWPCJogvOQkenaGwOreN3us3ZXddjfFK7I1EDsa5onWkPX1iyvUVejh
6vCvC0fOya95Kft5jH/BvuR48hGnatwsWYb8TPkindFYcwW1BdP/v3Me0rayNSopUWrFTU1b/mBz
tOx3Mpt2qlqcRBgr/03uzvmFGq7qjFqTx2uSxHF/UY5z+VRE8yMWyI9dx9PG5n/wz1GiXPkXZRqs
fjeyEpkWCUAMkzf1RxkjFbM8qqLNkiYgtPMeIUUhO1kaqK/MpNQNoFNkMBMcJR/mcjznCIc8XyO6
vYwd0twike1q5WzLYLyX9aOwtPAu32ahrQ+4PxtaUibr3sEKSO9Eu+jhRl/6+/+Ku2hSlWC6JWJP
dquTyRjrQwVdb4lHXSTUQCC3AvpoDdQTzp6heGrxTIH/DvR4U9GnX3hA3e5XDivI6sZ6l/gCbhrY
zXAZ3NlPKozwAkJeNuGvKuY+OP5GJCTrCKjkiurrEGvVuIRpYA7Ld/EVXIR2uD/1an4lWaKV3g1G
Pv/5V3jpV5jGQM/SbNKWJQPZQ/6BPSV1J6aYW65ieiKBN001hlmJ3gbhQPqc7mv51NKXWB8UGLk9
b2iyj4qPMjJXhtmXvKA+ANyQvJGJtmPS7/KS+Uh8IR3dFoOEIrUT1SFqAfX7Qf3CkDcvsGLm8vqj
cMURju9QE9msdqYpOCdjh61PH7D2JY9+EQNc+MDMIHCLQnnJZaxTpXO55dHLKTGciYm26AVKPaYH
14NxTaWWuBPnILI+LAEouPawXIat+VKfyY6wy+7LT8WaBFvCPl+QOtxtxwj1wauxDpf7FatQ+blC
q6Vrzn6j1bRgk04GcL8Qd7a/V+XlmW+8M+Y1rQ9nHDHDcI/3gAbSO1clVJqq0jWzGYZp2R3Ezqc5
Jxvzmkb7r8VKxnRHPIzqf3ZtnBAl68mxpFNoU/7nAxRuJ5j5eGeb0E2Tzd5NX5xFq3w66+PQLplA
MeoV5H+GsFlysEw3jdsNByETOt71fFCun8BuXpzd/c0+DdS3BsjhkDQKKi296E137MBMlPPHx7HN
ivdfqV0+d+5r52FdNGo/NJH/RmVjqsVduNVWVo5okOAiSoMAX9Pjjpxp4LSd+otiaOQhnvYZOvFt
5GES6K5hOF+RHgKU5PnhtgK6GmHsJy0PNPZxAaxHvw3gpN0IZcO6lyxfmlbjrh9hBU2WN6dAVlSU
2MQOBDI7JrAONHeh9QSVAg/HPh08NdeDTWUZ6p+qg+jXTf1V4GyL4n3MuLZ9MPoOlbryZ5w18kLw
udLGq4MrtOFlcP91jIzG6Nugk6L5lu14BWQ1i35mvcks2k62sFePKGHKJqywA3VWDV7Y0RZ1+zhe
m8gzXlgnJFQ/Njaa8r0qiM3maLVVWasVQ2qlbhsMnkoC8N7wr9NUx0Sa6MGFOJHXvhX1rKekmdo8
dDfVoI1M3nLuIhtTh3AOk8iL7o6vaCVMGk89Ju+SGF0qRn5E/YpwOr/kptVf5cs9Xi+AQxYxWbtm
iGbiykD8pBhcxc7alLI3uVUfyi6tnqWGY9conGYzsOKUhgzN/XpA9hh0PaA6SPdijKI179VD/334
5H+z2lZUFm/TPRRpboIdL4dC6l/ce2C3Ep/eKQDMPW4z1Dsg7jxh7me7aEuJTlUojqqUydzKoeqp
U3R7FmdzVnBTAfmsI7ifdJeVvBXQnc40VP9z1kFQu5r1Ep/gyu68m/hZgSoAnTffs/F3JeVDBHkv
NiKUwrRCtnOMHtBP98OIfFUWwEXl4hdLiDrpivkrOStmrh9LCdwZj9tsHDX30c+M/GhKNVYnsYKi
2XapgRuzmGGuCpMdBoiUFNhZQcqFezUI84wzFobJgsyywsOfYpLyxedANH8gx6mrcTaOkEjuCgXG
cy+agS0j2WN4DL9jIfl8uPbEsweymN5MfCmz2u4cwdcnfTt3gFnQ4gRBauuJTxJ05rVT+44o1mHw
tIHhGTx46OaWzHjdPMnu9R9Bfas49slHdvsmhaZjtKDINVc1Kv/QrgBrqAUAJW0wAMKSkh6filpf
zCXpy9IORPF3HDqJyAETdCn15PD/yeGvl4WfmIqGoKh861qzlErVIWQucZJzV3I9dqIF+DnZPNju
3ZKSOy76T1KOLDO9Dyy+mCWQr8T8N7gRrJkCxHoaqdfHG6l0Y28wSVRsyfhH4sQep0X3wT83KTtG
vLEr5LzB3umE4UrY3mx2va0KZff4rhzUwglIWHJ+KsMeOsy8dPBGm254sNtOKlQ1lYu4EaDduVwd
eY2Qo5MIi+uTDeJQd7WoIWdbBcInnfnL1b3EZjNun91rZgNuDqITTpEEZSDmnO6VqEO6eS8a0d8W
wgA0j/darsPTODLUPmQSHg+yNniIJWx2iX4gyJ524o5DSg6zMFUfvPjLUh0gD2pw3isxLPkvqN34
1RXSDwMg+v4ptsPRD6AlHD3pCXnAGfo92TgP1cd1OV7tZZicT4zvABpU2r798bKrnC7m9tryYX5y
1Rg308g/c3f1zhh+IDGp1KLZLd0Xr4SemscJaHl36qmbe7Pu4RB+SbxFhMof0PriXUIk5zRfWouC
iz7Loy/bHLOLE/MTktRad3ZJsWWNBFH9832TcM+6xoCzvZyai+TiswHvQN6uvj70ldzaO96f5r7P
8+Kk/3d1r6Ga8UtkEVXZ7BDbpWrPkFaLTMt/CoakDDkcUgVpQigOD7CAhtLQ7tdlLrOu38RPFe7L
i6J2L4zEnql4eP3oVeX3kMjE/8L2pdnB/nY2XsIohNt3bDuQrurEq2oRuASxw11S4la0ApBg+kJ/
Sz7sPTvESeSAFELSqJi+aQDidPgv3xcxILh23jSzeq0CZTMoR8lTWsP2g947heWaP0IVHV1u+CiK
WOwSbNgiTQrgpSchBe56hK78CuxmfcxTPhaEek8JjF5XMEXWfbN5bBAfUqG7ug48j1EjHxhjqdYR
6I05ZG+M4fVqSdPrGnZPLaOE1Jp023R1Ck1WzAnePanLRiYvEfvG5OfuzqL5pLRWKRzRFhi6mHEx
gIjSLD90gCCpoRiMaprN1N6DlKCG24tFAxsZj39715N/T7TWaCPh0D5hs/0nCpDZoL0wbU7QVwJF
uZZQ11vJlYKwCDdgXp154wAWwP1Fr7OT4knUsQVTsBL03gZzBv5sw3wpkk2W8lLd56KK5NT/AW8q
dRhZusfSjjLvOzHJ7NFtyj+jummh4I9xkfDw7oChpmhj+fi5muvd9LM+QkYgRAxyiJTxWzdAoYTh
zvb1KBvlh9He5APCXoYE+e99v+tbvHiCMztvvloO61kAzV1r3VH4SNjB3CYt+jwPXoo8XYWyQe1y
RiBe7Wam+uxEXeHeqnqJUDg2GrFtNJmuKNpKPnXm7aT1KSXOHoK45KiimQUzQgMIBOp73qYc0s2j
1y5M8DyPoDLaieAT/1T3PjRpipALDUS88hPF8rHf7iYbyH3xNFQwWClweoxwFCacXi4ItycMU6ZQ
6M0lvOuSAIHlv89yZSNskM2TbcSAZYFE5AQl8u4KK0XQ6xuwt0zje+oDNk9gV6wJgTZLI1pI21+i
Gtddf8ipAIQVSZirv1iuS4VT84C2nJ5sc/iZZYF6MWT3836W9BMM3+Z7HOKv7vauoQftUxrXXwHh
OLQ7BSO8cKsQp/wZl7GZSf7JOqNUwfoZn7kji9PR4eCaWv93Qf+58clVsjZdf/h2pW51MbIQx8E0
x9bRTLmhbe472mGk1QcC1pvZrP/zemP075JuFh1TbcCDezOgdk9Jmaw8BCDSLevGX6zEY90DgZzx
dmwSposipI7UYSVKOq0ctcBFmyQLk5wk7lin/0iIdw/6xvh8oG0sX8wyb5LKVht8TKWWZOeIF1m9
xRPZaC7b4N5HS9HghUDOw0L85bXiNm6YMiudnyVFj93xzXK2Y4mUSsmealxzHtI1e4xEhVWdWRQf
ujA0e9y3C56vreTbIZgpZh6AwxxhKeA9w7MMi4/GIjDt/5on09g5VTVoGUASt+LA/EMJzebA0fUW
0SLjVdkFkrgX9YTQga9cmvgCPNnnlnhlHAi/MfYTgjB6PQWqSyHJ2FilKJTnoY6A3k2gtMk/zLz4
48SZMC8/RT17vicAXxAbV69IIStaFSSYONonwvjnKmUzAA4NS3/fZjDDqFWu21k2as6ler55F8Yg
/y+VC6xD0pv8//9MIHzYUZFD7S5PuxW8GPVHHAhS2u8OiaLLesoNu8nsf4iYY7UIdIZ2xv4k7oRn
Cdp6Scm7+7uE0tfN8O8so24uB7Yasnbrn/cRmBqSqIvSiJ9LZCD32TPTCSzNqNQFztcjhbD1QlSS
SOmR5YVk/I45gJNq1zGj4u6D4yd/AQNxHRBjpa3T0u68rMXljvFY2EJfuISoYotjntcgHv3tTaZI
3YAKD8I3MLeNGlF9KU3kIp6WzDy23G8V+i/LWhdx2eeU/WfxWtHs9kK7MUZIu3MfVfiD/YaXlEq1
Vam0KCuN+LD/Hzl+mYKP5sp2wXnKX418/U1dKlSrUN4EUQ6ZdneNACm3jU+JWFCNSsGJpvxfH3zD
qMivGGGebPHgyHq1dE3nY34/lCsZrcLAt0Pwq7Ob7sQy1+fJyVcV2/1qod4F+qMvW1XiqLDLQamf
rUBSiK0EwsGd6fMekxCHeS/nuzOmsxJOeYF5sHafe2r+ViA8bLZyImBkya4z+cauc1avXiY1v4DZ
KyDZ/J4tbMnPF7LPiqHr3fFdy8IfLhpsdMHV9Qn9Ngi7X+2iax4U+BLFphiyTjXhsgP6cIk4d02I
2cSdhFHXAoN93c841k74cyd9JeXLSH9YFCxG7dYBpuzqGFQobe73tPCQABaoZBVIhITKtor4vzmX
lLlE/6DlbuMffYOlQS4TH5GYSc7Lpkba1viwL4IO4X11qwQSwL6+Cp9uKOQqOyTaolOUmsf1ApoQ
kaLf0pZhDHc0q/GsJTsVW/PawggwqK7YpeR7qGYlwtcLMGHtN+g8OMZ7aq89QjKl34alWLoGa6AV
H5YFMjd/StjzIOXESppEhbu8G3MC7RnAdRLoG9fD9fqjE2UdLxyoIDG0XG9IGYWnO3tfn5BnQx1M
PZGLmXSH2XBhEOoC+BTNBUvg86fpeYyo/oyLUXkxDSMj/PDYBRxo3XIIQ+eHQizEyAOcrKKgXB1V
wrI5pfQPHv1N+/4DCc7udvPgJA57JM6XDw+k+g6rjD8CsA8nbPA4gvjbm8FIpBEpsYQnw341SmAI
AYIlQocVdwpI8L9K8EgKHC1EqrgpiFPIeHRnULTc0tK9CsDeO4nn/72YbMxQ7S9B7IQuoUv8yuXT
Jw/LtivBrGhMdbal4LUw/Pmk2oq+d0Y5TpFi75ekc1VaEHM7yeluFGXeT3oyPc6ZND6bYLcJ8z3p
LHYf0SKpvfyoikHf2Wed/ErD/d4RICaz/I5E/LpAoWxFUtumUiMqgo9cNEKeK+tats+3P9Y5whn1
MQLBEfrCZwWsTqAhjBvTvl2iTRkMbbiMCdndrwQ8G9vV1zakQoAmYjOrJCIP79qh9EBb8CskoVxF
QyGoSeEPZ+TWnY7bX52ZKZk0Y86+ljSEtq5Y8BckvzsmOUtxxX4DFbAKszs9Lmlu7BIkbE78CeKH
iuEsHJdYt9tMY7ynxhb3FUPRrs3EALPFjCHnXJZLuOHw4rB6QJzzcS8ufzHmrRmjRmmqEoHmyTTt
06xjhAVlA3847acpJAPNpgF/YHMSMtaCztxRI7FffG96cQHhPSDD0ZnEx9V2VwQwfVEALr4mS2sJ
33898VQnaft9D9uYeFDp87Uo/Y29VBEMXnhzpmjUPZ6jpLYEHXy5o6pbw+lrumWzlS5+CfXaqk2z
/Wl/7ALfZsTQLzjXe4jxGTgabYZK1USC1B+ae70+UWR7OBGdWvU3/XqGrflsQXclran3D5xwyhfg
AOTy537EJqMJAYMSBMS+XmPR+eNUJ4J3v+Gnv0ql4yzhsmcHYUjUPVxcOoYVRMu5eXXa3O2/U6dx
bfDmm08U5K1mKBK7IuQYSJUboY8nwkNhbmw7hJewjmGx2kNxO8aQNvpgmR8dwoAUxxx71PEds/MM
XLvrJVHS1YlssDxAGix1APfZDZMAZpJHBVF9weuLdntRVAtAkpGAz4ug6rWnLv+8VjXphilE+Zjw
X0FUr/V0arrhlkqp2kmvSzZBQNMrx2FayCWBRYMW0rLkNddTJ5aE0zY991Al1zkPRvBDU/PwJXqC
sUwFbo37aydyO0PUlWLJ/OdqzsCHf4gaExeZ6sgoTJ+UXaVAAtRr8zLO7DW23lgazu1eIZEwA8Y1
Gd0illNeNQcGmxb7Z8xx6YsF77A30/uuQGm8oIh2n0TKnYvkzP0GCKyfNcti65Oy/sDJR+kKihE/
zzq3sftY1mmIiXkgOKHDjF5gSaCuK+lNOIllr3asmszGvpj6tnVaEHguO0idXG1ZQ1fgOGSlZ+P5
cMdoICwD3S5XDUPJ5+tIjIezNyCcS5HmPfl+pJKfijoCnXbms5QuEgdiebYEK/2f2aYtQ3X+V1lC
syMqeZYYjS8LXjZUUiOsNYLShMFQeA4ar/8OKJUIY++LKw7yOncNpQhANfUYkyaX42SNUl83Y0uQ
nhCeNVSDGwM55IgNmZtrFZ2G/26fLWlwuafRz7KS8OVBHaq5Zz18JEnjICtbLYazT/7ljQZEzonW
bCS5SSKeCBM7ySrrOlA7pSqgRbrCHo7fW93J6F7w67Pn+mtQxKSa/ynmKSO8ZhYIcUfvxbeYWAke
v+0kbZXuXj3h3kEXlUdMznKRR32RZK/4dgB7BDhAv2gBM1vDSWMtVFYXV660xNDPa6wpMM2oc9Uz
HhbDr7jLIiRAit8HqoDJK2wUV/K9JkSGnOe4wbmeddPk3zcV1HHolK8rnGh+FoOVIk/d2o62XVeS
yHKXF0NgKIovhrpHJA03HZw9BpgSUHnqSjaxOOH6fBdXFEphuQ/mdcem1cDKdXqpgPxZol47kleE
Fvy3y1A2c0g3mjeQ7PVUkYlR6XDQG06Iatze4F9z+EctlJ3V2a1iZJYNb0Z3y8+pBKqC09WWrSdD
lF+Mq6NcCLUkw09QFnnFGROOH5YZ1ov8IvGkgCEacgf3gZQbSqrEqQddD470rStgmq6rRLDPeL9T
hLpy57Tpq8zRl+VX9rcw5EqEb3+OPcPbyXTfgek048iSIDlnQcQ1EcqD/l5qUXAj+th2tz5LZAJo
6v2OVuXvNSFF72FjuxqLh84cLsMpllIkOeq+cCyVGQubqZcq32Zr71pZ3cS8CjTD3N7netMNdgCp
+58RJCzFWxJCdrAgPSC06V23/U8qoHLqrQuoHRuG8AfGD75gBB0+sy4//KwYopJLQalFCusN766c
TYyuIxRZY/hst9Pj7kC5CzoOTeggOC6BCvEdgf8z/4hWvUP4vydtYTUzZDXxsBn3GGdmsmNCqxl0
3UcOVY47wrIIjc0nHmFtXF0Y4BBVO4oD1TUPEYSo1wE4GSa+4GCedutOuLwRRoWZZVXpv4he0UsQ
NXGu6tPRcj6whS2rDF5dZSMF0DxApvGpCuoaDrLhlCmizU5YgVjcLBBg59LWEKnHCwHNid6gGuJI
S0MGjDlY34ULIPK3RKWZmlhbW2lPTNr+oCPyvkqIbkEuji7hR2R4aVnPjB8M14X2iSsumGKsj2JY
whNQV+lOLuRzFO/YMZOn/audO+7B8gbsUHCPCRvoViY6Sz2NslPcM6/IZQs8PiSsytY+Z8Ea48pm
XQ2MnYDIDSA2iRTRwdL+dYPTXwKGwBSjTv87tz4i31Dk+OWtVgqRZEoYB/3cKaMyKjJpINuBSxH1
gZzNU67+urEGjxfEiroIWIbR4C3xFNwJFrUHGYAIIj/SGfOkRdIpb34uoK/puMsClQDu9CJspepc
8fm2igX/mG8TIhPjh84KDEORCZCisfhTVzVpskdJ8bHBdZF60Nsf6yZO5E/sOGI11UNYV0zIzNe+
bg/W4Kk3F1lI2br75TGy6tWubn6dMqR8K3QgSjZQJ1S2bkNzfqo8pWjjf1wKOW6ZLwmv5C/IRDSc
OMJl65UQnlKaB5Q0ZEztp+yIz1QD8p1G3uBo3YUUlufdBmy0vOQBw7iOjlJyf3nkLtozXpiWhKIY
UADnUjCvEPuD6pJByTnoePFTeruhYMwTXOcDvMq1Tuu8Le0IEUZ65heuGGbwLRI8aL2Oekx84482
ZIzVVHbPrzW2lbowLR9bVGLJBqBc6O20PcSLVKX3LkHk9B7/tOwbG8H7ZOCA6/EWSfX0HZMz+V9C
3J/UtmhWpih62waOa+enCysxpriMHN+iSPfbIDDx368eM9ZxzQ9f053LC5z1QigqocMkVvxXpYWk
a5oZwy9uMvgg5hU8APy1VNRriMnfVhpCY7UXNCbBhEjvk/SjhonCg7szcQCNh9uHRizHB+eGhlIU
1PnfSRM85BhAPEwwHQkaD2DAeQac8ZB8o1vMxmujNqLIllpW61SWxRhi8Fe81Jm+kAS5ZP/aAkIK
PecApoA9sGplbPwKvWjtg+AoLlt8+m7SZgSxoGytx8JitOjYTQurcXgY1Q/vPxDkCepTcBcwLy86
OvH+qmj2+7LinCCfB2bIIO1570Z6M+S7kbck3p6B5ndpW02fHyNv5yBthy7RKG104VmY06kooR38
jIJUyoJxGohch7g7ZOO/gQ3YBuFIapRJzudc1ibvVlE/pf5kMrocjPWO8sbsa4NV6tv5KPUoDxg0
j3jD2xFDrCkEeRHtGcfkTfse97tSWlj5bXJlTsL3dFKfAfd+Ip47bSjeCNNZYml4vIUOv819mlQO
yDP0gtL8O5DQV3MUi2IPTl00iFGHzYgo6cPaFsgs5yFZZ1gsbQx9CxdhP7q5Df8zTCwImU+2evhf
t118m4l+Y38tAExRvhqUd1fMiMoN1311DgvjEjBUjCNZb6fpkolgzukEMclnpAIHCnvCvUnJr4uR
MNx7c5KwvB41mHgXdz2AzYYH97ZTUdDn66rwIZpEuWRn+eanGC65kgpjz9nAN9vfhXDKCg4D7XjR
Q9PkEkv91aHBzo3KtJU9SKjJnj6GBSI0E0Gvr5MhsFd4ZoYUnrpUpPpz/xNy/LQidswaVNNbiTfq
r4zUFLmi4sWOLkiX1LmKmSGnBDu41FxrUiuH5ldAUfppnJiDxuPy6MbjurScXTHosii9BAE0tk19
XlQxKHMvVhnDwmPZ1iZRz+bc1501MElbxKfCBKjJJ1rx7+bsCJJ9EmdDHZwEM72TrR9npDu5Wxll
wexQ7D+cFU8Vvq5iwnJS/xl55kJqyFN+I5cFBKrfMUbn/b0Av4VX4hcbfw/vIMH2hDxn8ncDJUbz
EPDdWUQCMcNTr79pQGdWxr+dqSHZ7oiJyMho5Og8eLim51zWuPc4hWggT7mgzCYqi+FO6T/IxNXl
0I+POs+MJh+oMVYlCnp1ASiJvuznsX0vj+6gne+uGFf9GQFprKdV5jd6vpnCk0d6a1beR+flg+bP
NbnDaFjVmSjeOv735O1k1UoMJatZVKHj6mGiGLAYfzEHU/gcA15uVTJrJZ1mF3O05dKT7fYc5pvs
E51PlyXkzU0TJY6jDhlAdshbKv3LXLIoOPHTs1Zpr1TLmnm92EzcqccER8tGCaj69dnGvUCkK7jQ
9j9a+vRjjVgdFwYEp+skL0CiQNZuplA1Od3gMhwv2FBFxACTeLGpGT0/extbpPnCDrJwoN5XKpHR
bXKaucyj9kuqWBRYqDvAStF5tyLVS6nvxXSSjY3oEl3VMWxas/I8q+NsqG+ZoO5eT/eI2XhQ13tS
87RyUH2sP6RVcYjf+gv9idNU/FXZjXXLkdj3oop5rkj9aovIWzvuXHUX34xHNJnNLfG2Gxt8THB7
0wO7XNkGnE42EeUTtOLWoiwxatgR0R6iFcXLNI+8aN2nP7pQyTyR97luEnz18RzeZ9ukBpYKNBHa
6khxUPjrb7dUKvOV1L6Vae7uI9yVJVsyJEKIUiWc1p47bkLxvkFTn5Sonl8nCAQTckAh0jwSBZLX
qdrCyzJfQQptgrP9rWZdXrBEcOVK9d0wqVx0iqimA6urkjefauax9nOTs092ShnGo1deoUmcOcKK
iZLm1ojPSTwW8vSxfrrdW9Bu3djHkC8f+C3g9cnKBJtpvYCWKUCwYLrhNsuUfzB+wEKHfkoymPVT
+dSSZp2NvpToNs5igCcT5uHuZjA/lWyPfDtmHHvarr7lza8HmVU0d9oYc0LJ4TabZ1sgf16tFDhR
ZyVbKQvVS+1+g/1/hQH2pCbLXGBGvSfCNEgSfk3CT2bIGodPzTmntK7rBZAeTHnszO6rIDXq8EMD
ZuhGKQ6DdJ0hL/25P+6yOPr8ygqYcm81UGLd9BajmiYGewLaMO7WU8oXF+PXgrXtRGrfTlGMgF/z
gElQZMYQFIwQnnA5N/nDwZAO8z5Up2BsZTjqEzVrAzHlgG2jXO7riPtwuL+CNvwOFsHgEAefpyiR
31eBwOVxm7RIug+KtGMEpvHX5Scj+N3GaVpaem/xgcA1vT9DKaPZ0kImp/6IDh8CMLJUPW+N1hsk
nozMUW9YXd7iVe0JHg+sPF81JhdhhO1Yd1q/C+CKOgGVGdDGNq9Tk1V45GiC+hbme5jfnRhtXlS3
LbMG+uZBLRwuEdqtBAL0uAfQ9HeduylikbHg4+2CCzGF6DSkMJYDUeUGoqoJyM/n2brEIeItOiKl
NdtUqDm9Xfxyb/X9gAJnGY70mNfZWQI6bBPOHLofbaRSy4R5F8i8UBlHzyi40ROuI/234H0WyDg8
DuRwT+k5UnK15s0PAt4uJzuIhFFDO5lp9sJCQ3cPm9o8RfdhOxXsCbQa2xy8nrFBNwIuvwGr427g
oLic6oHuDwLvmSiaB7SSO2oX62hOSudq/sMezwgCbReXY0ak4dyF0CiJQjVGx3aTZVbnW4FUSIbB
gUYiftMZ7wg7TlRO6GA8yARACPNQOw3MRxwHZqX80s9kHlSSkIUGvDwdwEvpdW/V/MBZFOtQEhW5
4Xy8hAgLkWQBHMdr0G36lDVOpw0ukbsHg6xQ4/AK7xHoT7n3Tetx+X+1yz+PB7AXkEiO4+PoN/qT
bM8YHD2gZ/O0NoqNS4/OjejAZ7KKlFjFnzfrzLcKYWuBaGzrYYXV2QHTRM2qkWvWB0sfnWTfjbzl
QY8d8v1Mm2ExLjnF0uM3HrU2z4fo3UrbNQDUGpkqJqoE1wmuGhw19ItpsEq+L2RStgs5+eU5py4X
06kLme0tXc8eU/MaRu4suvzLAMgrQJVD6qZFm5kgHdbH+nJyJWJomuQs8XGJhwd2ngBieRLDpNFR
v8GfqdJKwQ4gWVmaVumtj4ZujhbUumM8NBFavt2inAUUhYKP2Cj85ni69Ko2bPnmLlpRTUWyaF5q
dVgDveowHKAr4Y+lrIMBbDG2Ksfk3cpg1JLyp64AUctMvNhvpYaWfnAGOYCELMRZmVMMyda+LO9c
HmwA7+0yp7hkAFIgrD3ERlY49qAyTr0v+wItzNuObPpoicuizOfWovXwVPmnbtHhustNdZOtKGqq
HcCMYY0Aq/YcSfo+shyoIzVh0al/M48sjrqY+ft4lYvxC415Wz8CAGpnk0v3X3kTpTypU+P1KNb6
RX0Ui8p7ufjjTYXbg2miFUi4W1Qcl80N8jWrb/dFZEZNmchSU39kkgF/DTRzJ/efjunaDC4t+WdB
LzWUm+JHSiGk/9aCUZQ08B8Q6NrRYLpDDVLtn8i0WVdoCo4yVqG0j09dmL1ywzzN5FOIvQfdlylP
9jAlzlxTVEvQvFsp7O1pfiOQuQKQHcgH0ARPg/4+dzXrtj+734Lyb44TOg6F6AmB4RmKFnMBCp7d
kSMdO3fgzRjwJ9eg/R78sXE6coF2bFhdaHnQJzYFj092ABYhjP8OXrkEGcOdDTrbSXnh4tnp9Tcm
xRuiInlOwZMv4r0xoe5quV6oEvI1RyGliAWwcRAhkgyl+Ymh7vtYlXFU+HQDb73wpADV4KIEtbUB
PnuHH95D7M1q3P2spca7s9KhAa9P9t4bj/z5VTb1FrrkPLZjzQ4A2dywZB9H2sKkqh+v5bQeFD57
/EoQppDNXDok0sHHv7XyHO1rrx4iOP6wP3oIEP7R41mwmqkMCAuBjMvARmtMfTQIhO3caSVEVj3v
Z7U8XBskeKo+k83IGRbIfV3/If5J1W/XUInYwLEmbQicJ8MuwUZO2fL88bJkljoa7F/uW4rnxIq4
3/9Wrw/Ze7hLIxye/bHZAVQFymlhlOvMQQWCIEzqgrwECkN+PBfcL5lwba2RpNg1wTQNGS0quW1n
xgbiwNyx4v6AKcuvwqnrAO5b4HmT0SXFxzkBSqKkizQPh8D9kpks2YJZ30CTHdzsuAY90iE3oLs8
g4iUbvMgmSRoWBgcBNLfIGvvi88eJYqUTuAGc5uofrpZ9/N9o4kHJ//63EXd+FyqEtai4QTrrHys
SzCpeHSPuDofVQX9WyM1QySZTElfoPTjR0uYPT1huPLF6w==
`protect end_protected
