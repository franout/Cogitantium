// Register NVDLA_MCIF_CFG_RD_WEIGHT_0_0
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0					32'h2000
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_BDMA_RANGE			7:0
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_BDMA_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_SDP_RANGE			15:8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_SDP_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_PDP_RANGE			23:16
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_PDP_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_CDP_RANGE			31:24
#define NVDLA_MCIF_CFG_RD_WEIGHT_0_0_RD_WEIGHT_CDP_SIZE				8


// Register NVDLA_MCIF_CFG_RD_WEIGHT_1_0
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0					32'h2004
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_B_RANGE			7:0
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_B_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_N_RANGE			15:8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_N_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_E_RANGE			23:16
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_SDP_E_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_CDMA_DAT_RANGE			31:24
#define NVDLA_MCIF_CFG_RD_WEIGHT_1_0_RD_WEIGHT_CDMA_DAT_SIZE				8


// Register NVDLA_MCIF_CFG_RD_WEIGHT_2_0
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0					32'h2008
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_CDMA_WT_RANGE			7:0
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_CDMA_WT_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RBK_RANGE			15:8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RBK_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_1_RANGE			23:16
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_1_SIZE				8
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_0_RANGE			31:24
#define NVDLA_MCIF_CFG_RD_WEIGHT_2_0_RD_WEIGHT_RSV_0_SIZE				8


// Register NVDLA_MCIF_CFG_WR_WEIGHT_0_0
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0					32'h200c
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_BDMA_RANGE			7:0
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_BDMA_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_SDP_RANGE			15:8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_SDP_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_PDP_RANGE			23:16
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_PDP_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_CDP_RANGE			31:24
#define NVDLA_MCIF_CFG_WR_WEIGHT_0_0_WR_WEIGHT_CDP_SIZE				8


// Register NVDLA_MCIF_CFG_WR_WEIGHT_1_0
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0					32'h2010
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RBK_RANGE			7:0
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RBK_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_2_RANGE			15:8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_2_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_1_RANGE			23:16
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_1_SIZE				8
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_0_RANGE			31:24
#define NVDLA_MCIF_CFG_WR_WEIGHT_1_0_WR_WEIGHT_RSV_0_SIZE				8


// Register NVDLA_MCIF_CFG_OUTSTANDING_CNT_0
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0					32'h2014
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_RD_OS_CNT_RANGE			7:0
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_RD_OS_CNT_SIZE				8
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_WR_OS_CNT_RANGE			15:8
#define NVDLA_MCIF_CFG_OUTSTANDING_CNT_0_WR_OS_CNT_SIZE				8


// Register NVDLA_MCIF_STATUS_0
#define NVDLA_MCIF_STATUS_0					32'h2018
#define NVDLA_MCIF_STATUS_0_IDLE_RANGE			8:8
#define NVDLA_MCIF_STATUS_0_IDLE_SIZE				1
#define NVDLA_MCIF_STATUS_0_IDLE_NO			1'h0
#define NVDLA_MCIF_STATUS_0_IDLE_YES			1'h1



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_MCIF	32'h2000
