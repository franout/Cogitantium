// Register NVDLA_CMAC_A_S_STATUS_0
#define NVDLA_CMAC_A_S_STATUS_0					32'h5000
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_RANGE			1:0
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_SIZE				2
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_IDLE			2'h0
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_RUNNING			2'h1
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_0_PENDING			2'h2
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_RANGE			17:16
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_SIZE				2
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_IDLE			2'h0
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_RUNNING			2'h1
#define NVDLA_CMAC_A_S_STATUS_0_STATUS_1_PENDING			2'h2


// Register NVDLA_CMAC_A_S_POINTER_0
#define NVDLA_CMAC_A_S_POINTER_0					32'h5004
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_RANGE			0:0
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_SIZE				1
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_GROUP_0			1'h0
#define NVDLA_CMAC_A_S_POINTER_0_PRODUCER_GROUP_1			1'h1
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_RANGE			16:16
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_SIZE				1
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_GROUP_0			1'h0
#define NVDLA_CMAC_A_S_POINTER_0_CONSUMER_GROUP_1			1'h1


// Register NVDLA_CMAC_A_D_OP_ENABLE_0
#define NVDLA_CMAC_A_D_OP_ENABLE_0					32'h5008
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_RANGE			0:0
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_SIZE				1
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_DISABLE			1'h0
#define NVDLA_CMAC_A_D_OP_ENABLE_0_OP_EN_ENABLE			1'h1


// Register NVDLA_CMAC_A_D_MISC_CFG_0
#define NVDLA_CMAC_A_D_MISC_CFG_0					32'h500c
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_RANGE			0:0
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_SIZE				1
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_DIRECT			1'h0
#define NVDLA_CMAC_A_D_MISC_CFG_0_CONV_MODE_WINOGRAD			1'h1
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_RANGE			13:12
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_SIZE				2
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_INT8			2'h0
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_INT16			2'h1
#define NVDLA_CMAC_A_D_MISC_CFG_0_PROC_PRECISION_FP16			2'h2



//
// ADDRESS SPACES
//

#define BASE_ADDRESS_NVDLA_CMAC_A	32'h5000
